magic
tech scmos
timestamp 1619549734
<< nwell >>
rect 0 0 24 48
rect 30 0 54 48
<< ntransistor >>
rect 11 -43 13 -8
rect 41 -43 43 -8
<< ptransistor >>
rect 11 12 13 17
rect 41 12 43 17
<< ndiffusion >>
rect 10 -43 11 -8
rect 13 -43 14 -8
rect 40 -43 41 -8
rect 43 -43 44 -8
<< pdiffusion >>
rect 10 12 11 17
rect 13 12 14 17
rect 40 12 41 17
rect 43 12 44 17
<< ndcontact >>
rect 6 -43 10 -8
rect 14 -43 18 -8
rect 36 -43 40 -8
rect 44 -43 48 -8
<< pdcontact >>
rect 6 12 10 17
rect 14 12 18 17
rect 36 12 40 17
rect 44 12 48 17
<< polysilicon >>
rect 11 17 13 22
rect 41 17 43 21
rect 11 -8 13 12
rect 41 -8 43 12
rect 11 -46 13 -43
rect 41 -46 43 -43
<< polycontact >>
rect 7 -5 11 -1
rect 37 -5 41 -1
<< metal1 >>
rect 0 48 54 51
rect 6 17 10 48
rect 36 17 40 48
rect 14 -1 18 12
rect 0 -5 7 -1
rect 14 -5 37 -1
rect 44 -2 48 12
rect 14 -8 18 -5
rect 44 -6 54 -2
rect 44 -8 48 -6
rect 6 -46 10 -43
rect 36 -46 40 -43
rect 0 -49 54 -46
<< end >>
