magic
tech scmos
timestamp 1619531845
<< metal1 >>
rect -124 168 -120 169
rect -107 168 -102 257
rect 125 223 129 261
rect 42 208 47 222
rect 131 179 136 185
rect -73 174 136 179
rect 228 178 233 187
rect 176 173 233 178
rect 326 177 331 185
rect 291 172 331 177
rect 341 168 345 170
rect -124 165 12 168
rect -124 -34 -120 165
rect 9 111 13 113
rect 56 111 60 113
rect 107 104 111 106
rect 152 104 156 106
rect 206 104 210 106
rect 252 104 256 106
rect 303 104 307 106
rect 350 104 354 106
rect 356 66 360 68
rect 136 -6 141 5
rect -100 -10 141 -6
rect 322 -52 327 -47
rect 322 -89 327 -57
rect 322 -93 334 -89
rect 378 -128 381 -58
rect -62 -215 -57 -179
rect -111 -262 50 -257
rect 303 -273 307 -224
rect 497 -273 563 -272
rect 390 -276 450 -273
rect 500 -275 563 -273
rect 558 -286 563 -275
rect 500 -330 562 -326
rect 43 -335 48 -330
rect 2 -373 9 -370
rect 427 -373 487 -370
rect 500 -373 565 -370
rect 112 -501 116 -497
rect 107 -505 117 -501
rect 215 -505 219 -497
rect 317 -501 321 -497
rect 416 -501 420 -497
rect 317 -505 320 -501
rect 418 -505 419 -501
rect 219 -548 224 -545
rect 320 -548 325 -545
rect 419 -548 424 -545
<< m2contact >>
rect 42 222 47 227
rect 137 211 142 216
rect 234 211 239 216
rect 377 63 382 68
rect 233 0 238 5
rect 331 -1 336 4
rect -105 -11 -100 -6
rect 322 -47 327 -42
rect -105 -84 -100 -79
rect 377 -58 382 -53
rect 555 -56 560 -51
rect -163 -184 -158 -179
rect -62 -220 -57 -215
rect 446 -330 451 -325
<< metal2 >>
rect -421 -618 -416 261
rect -251 247 -246 252
rect 277 249 282 250
rect 548 236 553 249
rect -180 222 42 227
rect -180 -95 -174 222
rect 94 212 137 216
rect 94 -4 97 212
rect 189 211 234 216
rect 131 174 136 182
rect -105 -71 -100 -11
rect -111 -72 -100 -71
rect -105 -79 -100 -72
rect -36 -10 97 -4
rect -36 -93 -31 -10
rect 189 -11 193 211
rect 176 -16 193 -11
rect 233 -25 238 0
rect 78 -28 238 -25
rect 322 -1 331 4
rect 78 -88 83 -28
rect 322 -42 327 -1
rect 377 -53 382 63
rect -163 -231 -158 -184
rect -57 -220 200 -216
rect -163 -236 105 -231
rect 100 -361 105 -236
rect 195 -361 200 -220
rect 555 -247 560 -56
rect 446 -251 560 -247
rect 446 -325 451 -251
rect 385 -434 504 -433
rect 385 -438 505 -434
rect 502 -596 505 -438
rect -421 -621 -277 -618
<< m3contact >>
rect -251 242 -246 247
rect 11 245 16 250
rect 277 244 282 249
rect 548 231 553 236
rect 36 147 41 152
rect -111 -71 -105 -66
rect 78 -146 83 -141
<< m123contact >>
rect -78 174 -73 179
rect -1 106 4 111
rect 38 0 43 5
rect 332 211 337 216
rect 171 173 176 178
rect 102 106 107 111
rect 286 172 291 177
rect 197 106 202 111
rect 295 106 300 111
rect 171 -16 176 -11
rect 322 -57 327 -52
rect 171 -92 176 -87
rect 505 -171 510 -166
rect -2 -180 3 -175
rect 227 -179 232 -174
rect -116 -262 -111 -257
rect 50 -262 55 -257
rect -2 -335 3 -330
rect 38 -335 43 -330
rect 142 -335 147 -330
rect 239 -335 244 -330
rect 293 -335 298 -330
rect 337 -335 342 -330
rect 117 -506 122 -501
rect 219 -506 224 -501
rect 320 -506 325 -501
rect 419 -506 424 -501
rect 256 -553 261 -548
<< metal3 >>
rect -246 242 -150 247
rect -154 111 -150 242
rect -141 152 -136 261
rect -129 179 -124 261
rect 16 245 107 249
rect -129 174 -78 179
rect -141 147 36 152
rect 102 111 107 245
rect 137 239 142 261
rect 392 252 397 261
rect 191 244 277 249
rect 286 247 397 252
rect 137 234 176 239
rect 171 178 176 234
rect -154 106 -1 111
rect 4 106 5 111
rect 191 111 196 244
rect 286 177 291 247
rect 296 235 548 236
rect 295 231 548 235
rect 295 111 300 231
rect 337 211 435 216
rect 191 106 197 111
rect -116 -257 -111 -66
rect 3 -180 4 -175
rect -2 -330 1 -180
rect 38 -330 42 0
rect 171 -87 176 -16
rect 327 -57 374 -52
rect 72 -146 78 -141
rect 72 -249 77 -146
rect 227 -240 232 -179
rect 369 -229 374 -57
rect 430 -166 435 211
rect 430 -171 505 -166
rect 337 -234 374 -229
rect 227 -244 298 -240
rect 72 -254 244 -249
rect 55 -262 147 -258
rect 142 -330 147 -262
rect 239 -330 244 -254
rect 293 -330 298 -244
rect 337 -330 342 -234
rect 117 -576 122 -506
rect -247 -581 122 -576
rect -247 -596 -242 -581
rect 219 -591 224 -506
rect 15 -596 224 -591
rect 256 -596 261 -553
rect 320 -554 325 -506
rect 281 -560 325 -554
rect 419 -554 424 -506
rect 419 -558 557 -554
rect 281 -596 287 -560
rect 552 -596 557 -558
use pg  pg_0
timestamp 1619531378
transform 1 0 9 0 1 68
box -9 -68 382 155
use cla  cla_0
timestamp 1619531378
transform 1 0 -171 0 1 -131
box -20 -95 741 100
use sum  sum_0
timestamp 1619527417
transform 1 0 7 0 1 -373
box -9 -175 424 100
use buff  buff_0
timestamp 1619185680
transform 1 0 446 0 1 -324
box 0 -49 54 51
use dff  dff_4
timestamp 1619465570
transform 1 0 581 0 1 -373
box 0 -201 239 89
<< labels >>
rlabel space 497 -328 497 -328 1 dc4
rlabel metal1 112 -501 116 -497 1 ds1
rlabel metal1 215 -501 219 -497 1 ds2
rlabel metal1 317 -501 321 -497 1 ds3
rlabel metal1 416 -501 420 -497 1 ds4
rlabel metal1 9 111 13 113 1 a1
rlabel metal1 56 111 60 113 1 b1
rlabel metal1 107 104 111 106 1 a2
rlabel metal1 152 104 156 106 1 b2
rlabel metal1 206 104 210 106 1 a3
rlabel metal1 252 104 256 106 1 b3
rlabel metal1 303 104 307 106 1 a4
rlabel metal1 350 104 354 106 1 b4
rlabel metal1 341 168 345 170 1 vdd
rlabel metal1 356 66 360 68 1 gnd
<< end >>
