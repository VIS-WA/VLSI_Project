magic
tech scmos
timestamp 1619527417
<< nwell >>
rect 95 50 119 74
rect 143 50 167 74
rect 192 50 216 74
rect 240 50 264 74
rect 290 50 314 74
rect 338 50 362 74
<< ntransistor >>
rect 106 15 108 20
rect 154 15 156 20
rect 203 15 205 20
rect 251 15 253 20
rect 301 15 303 20
rect 349 15 351 20
<< ptransistor >>
rect 106 58 108 68
rect 154 58 156 68
rect 203 58 205 68
rect 251 58 253 68
rect 301 58 303 68
rect 349 58 351 68
<< ndiffusion >>
rect 105 15 106 20
rect 108 15 109 20
rect 153 15 154 20
rect 156 15 157 20
rect 202 15 203 20
rect 205 15 206 20
rect 250 15 251 20
rect 253 15 254 20
rect 300 15 301 20
rect 303 15 304 20
rect 348 15 349 20
rect 351 15 352 20
<< pdiffusion >>
rect 105 58 106 68
rect 108 58 109 68
rect 153 58 154 68
rect 156 58 157 68
rect 202 58 203 68
rect 205 58 206 68
rect 250 58 251 68
rect 253 58 254 68
rect 300 58 301 68
rect 303 58 304 68
rect 348 58 349 68
rect 351 58 352 68
<< ndcontact >>
rect 101 15 105 20
rect 109 15 113 20
rect 149 15 153 20
rect 157 15 161 20
rect 198 15 202 20
rect 206 15 210 20
rect 246 15 250 20
rect 254 15 258 20
rect 296 15 300 20
rect 304 15 308 20
rect 344 15 348 20
rect 352 15 356 20
<< pdcontact >>
rect 101 58 105 68
rect 109 58 113 68
rect 149 58 153 68
rect 157 58 161 68
rect 198 58 202 68
rect 206 58 210 68
rect 246 58 250 68
rect 254 58 258 68
rect 296 58 300 68
rect 304 58 308 68
rect 344 58 348 68
rect 352 58 356 68
<< polysilicon >>
rect 106 68 108 71
rect 154 68 156 71
rect 203 68 205 71
rect 251 68 253 71
rect 301 68 303 71
rect 349 68 351 71
rect 106 20 108 58
rect 154 20 156 58
rect 203 20 205 58
rect 251 20 253 58
rect 301 20 303 58
rect 349 20 351 58
rect 106 12 108 15
rect 154 12 156 15
rect 203 12 205 15
rect 251 12 253 15
rect 301 12 303 15
rect 349 12 351 15
<< polycontact >>
rect 101 38 106 43
rect 149 38 154 43
rect 198 38 203 43
rect 246 38 251 43
rect 296 38 301 43
rect 344 38 349 43
<< metal1 >>
rect 24 97 378 100
rect 101 68 105 97
rect 149 68 153 97
rect 198 68 202 97
rect 246 68 250 97
rect 296 68 300 97
rect 344 68 348 97
rect -9 38 0 43
rect 37 38 48 43
rect 93 38 101 43
rect -9 -44 -4 38
rect 24 26 28 31
rect 37 13 42 38
rect 72 26 74 31
rect 93 17 98 38
rect 109 31 113 58
rect 135 38 149 43
rect 109 26 119 31
rect 109 20 113 26
rect 135 17 140 38
rect 157 31 161 58
rect 188 38 198 43
rect 157 26 169 31
rect 157 20 161 26
rect 101 3 105 15
rect 188 17 193 38
rect 206 31 210 58
rect 232 38 246 43
rect 206 26 216 31
rect 206 20 210 26
rect 149 3 153 15
rect 232 17 237 38
rect 254 31 258 58
rect 286 38 296 43
rect 254 26 266 31
rect 254 20 258 26
rect 198 3 202 15
rect 286 17 291 38
rect 304 31 308 58
rect 330 38 344 43
rect 304 26 314 31
rect 304 20 308 26
rect 246 3 250 15
rect 330 17 335 38
rect 352 31 356 58
rect 352 26 364 31
rect 352 20 356 26
rect 296 3 300 15
rect 344 3 348 15
rect 24 0 424 3
rect 20 -44 25 -29
rect 37 -44 42 -9
rect 52 -44 57 -18
rect 93 -39 98 -8
rect 118 -39 123 -29
rect 135 -39 140 -8
rect 150 -39 155 -17
rect 188 -39 193 -8
rect 215 -39 220 -29
rect 232 -39 237 -8
rect 247 -39 252 -17
rect 286 -39 291 -8
rect 93 -44 106 -39
rect 188 -44 204 -39
rect 286 -40 303 -39
rect 313 -40 318 -29
rect 330 -40 335 -8
rect 345 -40 350 -17
rect 286 -44 302 -40
rect -9 -50 8 -44
rect 29 -128 34 -68
rect 100 -78 415 -75
rect 29 -132 46 -128
rect 420 -172 424 0
rect 100 -175 424 -172
<< m2contact >>
rect 378 95 383 100
rect 28 26 33 31
rect 69 21 74 26
rect 37 8 42 13
rect 119 26 124 31
rect 93 12 98 17
rect 164 21 169 26
rect 135 12 140 17
rect 216 26 221 31
rect 188 12 193 17
rect 261 21 266 26
rect 232 12 237 17
rect 314 26 319 31
rect 286 12 291 17
rect 359 21 364 26
rect 330 12 335 17
rect 37 -9 42 -4
rect 20 -29 25 -23
rect 93 -8 98 -3
rect 52 -18 57 -13
rect 135 -8 140 -3
rect 118 -29 123 -23
rect 188 -8 193 -3
rect 150 -17 155 -12
rect 232 -8 237 -3
rect 215 -29 220 -23
rect 286 -8 291 -3
rect 247 -17 252 -12
rect 330 -8 335 -3
rect 313 -29 318 -23
rect 345 -17 350 -12
rect 127 -68 132 -63
rect 224 -68 229 -63
rect 322 -69 327 -64
rect 378 -75 383 -70
rect 149 -132 154 -127
rect 251 -132 256 -127
rect 352 -132 357 -127
<< metal2 >>
rect 28 -13 33 26
rect 37 -4 42 8
rect 28 -18 52 -13
rect 69 -23 74 21
rect 93 -3 98 12
rect 119 -12 124 26
rect 135 -3 140 12
rect 119 -17 150 -12
rect 164 -23 169 21
rect 188 -3 193 12
rect 216 -12 221 26
rect 232 -3 237 12
rect 216 -17 247 -12
rect 261 -23 266 21
rect 286 -3 291 12
rect 314 -12 319 26
rect 330 -3 335 12
rect 314 -17 345 -12
rect 359 -23 364 21
rect 25 -29 74 -23
rect 123 -29 169 -23
rect 220 -29 266 -23
rect 318 -29 364 -23
rect 127 -128 132 -68
rect 127 -132 149 -128
rect 224 -128 229 -68
rect 224 -132 251 -128
rect 322 -128 327 -69
rect 378 -70 383 95
rect 322 -132 352 -128
use not  not_0
timestamp 1619185627
transform 1 0 0 0 1 47
box 0 -47 24 53
use not  not_1
timestamp 1619185627
transform 1 0 48 0 1 47
box 0 -47 24 53
use xor  xor_0
timestamp 1618556316
transform 0 -1 32 1 0 -68
box 0 -28 24 30
use xor  xor_1
timestamp 1618556316
transform 0 -1 130 1 0 -63
box 0 -28 24 30
use xor  xor_2
timestamp 1618556316
transform 0 -1 227 1 0 -63
box 0 -28 24 30
use xor  xor_3
timestamp 1618556316
transform 0 -1 325 1 0 -64
box 0 -28 24 30
use buff  buff_0
timestamp 1619185680
transform 1 0 46 0 1 -126
box 0 -49 54 51
use buff  buff_1
timestamp 1619185680
transform 1 0 154 0 1 -126
box 0 -49 54 51
use buff  buff_2
timestamp 1619185680
transform 1 0 256 0 1 -126
box 0 -49 54 51
use buff  buff_3
timestamp 1619185680
transform 1 0 357 0 1 -126
box 0 -49 54 51
<< labels >>
rlabel metal1 347 1 347 1 1 gnd
rlabel metal1 343 99 343 99 4 vdd
rlabel metal1 -4 40 -4 40 3 c0
rlabel space 18 28 18 28 1 c0_b
rlabel metal1 45 41 45 41 1 p1
rlabel space 70 28 70 28 1 p1_b
rlabel metal1 98 40 98 40 1 c1
rlabel metal1 116 29 116 29 1 c1_b
rlabel metal1 143 41 143 41 1 p2
rlabel metal1 166 28 166 28 1 p2_b
rlabel metal1 193 41 193 41 1 c2
rlabel metal1 213 28 213 28 1 c2_b
rlabel metal1 239 41 239 41 1 p3
rlabel metal1 261 29 261 29 1 p3_b
rlabel metal1 293 41 293 41 1 c3
rlabel metal1 311 29 311 29 1 c3_b
rlabel metal1 340 41 340 41 1 p4
rlabel metal1 360 29 360 29 7 p4_b
rlabel space 31 -60 31 -60 1 ss1
rlabel space 130 -56 130 -56 1 ss2
rlabel space 227 -56 227 -56 1 ss3
rlabel space 325 -57 325 -57 1 ss4
<< end >>
