magic
tech scmos
timestamp 1613729823
<< nwell >>
rect -8 -5 17 40
<< ntransistor >>
rect 4 -23 6 -13
<< ptransistor >>
rect 4 1 6 26
<< ndiffusion >>
rect 3 -23 4 -13
rect 6 -23 7 -13
<< pdiffusion >>
rect 3 1 4 26
rect 6 1 7 26
<< ndcontact >>
rect -1 -23 3 -13
rect 7 -23 11 -13
<< pdcontact >>
rect -1 1 3 26
rect 7 1 11 26
<< polysilicon >>
rect 4 26 6 29
rect 4 -13 6 1
rect 4 -26 6 -23
<< polycontact >>
rect 0 -10 4 -6
<< metal1 >>
rect -8 36 17 40
rect -1 26 3 36
rect 7 -6 11 1
rect -11 -10 0 -6
rect 7 -10 20 -6
rect 7 -13 11 -10
rect -1 -33 3 -23
rect -8 -37 17 -33
<< labels >>
rlabel metal1 -8 -8 -8 -8 3 in
rlabel metal1 19 -8 19 -8 7 out
rlabel metal1 16 39 16 39 6 vdd
rlabel metal1 16 -35 16 -35 8 gnd
<< end >>
