4 bit CLA
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={5*LAMBDA}
.param width_P={10*LAMBDA}
.global gnd vdd

Vdd vdd gnd 'SUPPLY'

.option scale=0.09u

va1 a 0 pulse 0 1.8 0ns 0ns 0ns 5ns 10ns
va2 b 0 pulse 0 1.8 0ns 0ns 0ns 10ns 20ns
va3 c 0 pulse 0 1.8 0ns 0ns 0ns 15ns 30ns


M1000 out b vdd vdd CMOSP w=10 l=2
+  ad=150 pd=90 as=150 ps=90
M1001 out c vdd vdd CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out a vdd vdd CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 x a y Gnd CMOSN w=5 l=2
+  ad=50 pd=40 as=50 ps=40
M1004 out b x Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1005 y c gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=25 ps=20
C0 x a 0.11fF
C1 c vdd 0.08fF
C2 a vdd 0.27fF
C3 out a 0.09fF
C4 c out 0.15fF
C5 vdd a 0.58fF
C6 out vdd 0.07fF
C7 a vdd 0.22fF
C8 x out 0.08fF
C9 vdd vdd 0.08fF
C10 b a 0.31fF
C11 out vdd 0.04fF
C12 vdd vdd 0.06fF
C13 out vdd 0.34fF
C14 x b 0.02fF
C15 out vdd 0.04fF
C16 b vdd 0.08fF
C17 out b 0.17fF
C18 vdd vdd 0.07fF
C19 gnd y 0.08fF
C20 y c 0.08fF
C21 c a 0.01fF
C22 y x 0.09fF


.tran 0.1n 40n

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7)
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7)


run
plot v(a) v(b)+2 v(c)+4 v(out)+6
.endc
