magic
tech scmos
timestamp 1619530824
<< nwell >>
rect -341 844 -317 873
rect -306 844 -282 873
rect -175 844 -151 873
rect -140 844 -116 873
rect -38 844 -14 873
rect -3 844 21 873
rect 128 844 152 873
rect 163 844 187 873
rect 258 844 282 873
rect 293 844 317 873
rect 424 844 448 873
rect 459 844 483 873
rect 570 844 594 873
rect 605 844 629 873
rect 736 844 760 873
rect 771 844 795 873
rect -341 666 -317 724
rect -306 666 -282 724
rect -271 666 -247 695
rect -175 666 -151 724
rect -140 666 -116 724
rect -38 666 -14 724
rect -3 666 21 724
rect 32 666 56 695
rect 128 666 152 724
rect 163 666 187 724
rect 258 666 282 724
rect 293 666 317 724
rect 328 666 352 695
rect 424 666 448 724
rect 459 666 483 724
rect 570 666 594 724
rect 605 666 629 724
rect 640 666 664 695
rect 736 666 760 724
rect 771 666 795 724
rect -290 -679 -266 -650
rect -255 -679 -231 -650
rect -124 -679 -100 -650
rect -89 -679 -65 -650
rect 13 -679 37 -650
rect 48 -679 72 -650
rect 179 -679 203 -650
rect 214 -679 238 -650
rect 309 -679 333 -650
rect 344 -679 368 -650
rect 475 -679 499 -650
rect 510 -679 534 -650
rect 621 -679 645 -650
rect 656 -679 680 -650
rect 787 -679 811 -650
rect 822 -679 846 -650
rect -290 -857 -266 -799
rect -255 -857 -231 -799
rect -220 -857 -196 -828
rect -124 -857 -100 -799
rect -89 -857 -65 -799
rect 13 -857 37 -799
rect 48 -857 72 -799
rect 83 -857 107 -828
rect 179 -857 203 -799
rect 214 -857 238 -799
rect 309 -857 333 -799
rect 344 -857 368 -799
rect 379 -857 403 -828
rect 475 -857 499 -799
rect 510 -857 534 -799
rect 621 -857 645 -799
rect 656 -857 680 -799
rect 691 -857 715 -828
rect 787 -857 811 -799
rect 822 -857 846 -799
<< ntransistor >>
rect -312 817 -310 822
rect -146 817 -144 822
rect -9 817 -7 822
rect 157 817 159 822
rect 287 817 289 822
rect 453 817 455 822
rect 599 817 601 822
rect 765 817 767 822
rect -312 797 -310 802
rect -146 797 -144 802
rect -9 797 -7 802
rect 157 797 159 802
rect 287 797 289 802
rect 453 797 455 802
rect 599 797 601 802
rect 765 797 767 802
rect -312 766 -310 771
rect -146 766 -144 771
rect -9 766 -7 771
rect 157 766 159 771
rect 287 766 289 771
rect 453 766 455 771
rect 599 766 601 771
rect 765 766 767 771
rect -312 746 -310 751
rect -146 746 -144 751
rect -9 746 -7 751
rect 157 746 159 751
rect 287 746 289 751
rect 453 746 455 751
rect 599 746 601 751
rect 765 746 767 751
rect -312 639 -310 644
rect -312 615 -310 620
rect -146 639 -144 644
rect -9 639 -7 644
rect -146 619 -144 624
rect -9 615 -7 620
rect 157 639 159 644
rect 287 639 289 644
rect 157 619 159 624
rect 287 615 289 620
rect 453 639 455 644
rect 599 639 601 644
rect 453 619 455 624
rect 599 615 601 620
rect 765 639 767 644
rect 765 619 767 624
rect -312 596 -310 601
rect -9 596 -7 601
rect 287 596 289 601
rect 599 596 601 601
rect -261 -706 -259 -701
rect -95 -706 -93 -701
rect 42 -706 44 -701
rect 208 -706 210 -701
rect 338 -706 340 -701
rect 504 -706 506 -701
rect 650 -706 652 -701
rect 816 -706 818 -701
rect -261 -726 -259 -721
rect -95 -726 -93 -721
rect 42 -726 44 -721
rect 208 -726 210 -721
rect 338 -726 340 -721
rect 504 -726 506 -721
rect 650 -726 652 -721
rect 816 -726 818 -721
rect -261 -757 -259 -752
rect -95 -757 -93 -752
rect 42 -757 44 -752
rect 208 -757 210 -752
rect 338 -757 340 -752
rect 504 -757 506 -752
rect 650 -757 652 -752
rect 816 -757 818 -752
rect -261 -777 -259 -772
rect -95 -777 -93 -772
rect 42 -777 44 -772
rect 208 -777 210 -772
rect 338 -777 340 -772
rect 504 -777 506 -772
rect 650 -777 652 -772
rect 816 -777 818 -772
rect -261 -884 -259 -879
rect -261 -908 -259 -903
rect -95 -884 -93 -879
rect 42 -884 44 -879
rect -95 -904 -93 -899
rect 42 -908 44 -903
rect 208 -884 210 -879
rect 338 -884 340 -879
rect 208 -904 210 -899
rect 338 -908 340 -903
rect 504 -884 506 -879
rect 650 -884 652 -879
rect 504 -904 506 -899
rect 650 -908 652 -903
rect 816 -884 818 -879
rect 816 -904 818 -899
rect -261 -927 -259 -922
rect 42 -927 44 -922
rect 338 -927 340 -922
rect 650 -927 652 -922
<< ptransistor >>
rect -330 852 -328 862
rect -295 852 -293 862
rect -164 852 -162 862
rect -129 852 -127 862
rect -27 852 -25 862
rect 8 852 10 862
rect 139 852 141 862
rect 174 852 176 862
rect 269 852 271 862
rect 304 852 306 862
rect 435 852 437 862
rect 470 852 472 862
rect 581 852 583 862
rect 616 852 618 862
rect 747 852 749 862
rect 782 852 784 862
rect -330 706 -328 716
rect -295 706 -293 716
rect -164 706 -162 716
rect -129 706 -127 716
rect -27 706 -25 716
rect 8 706 10 716
rect 139 706 141 716
rect 174 706 176 716
rect 269 706 271 716
rect 304 706 306 716
rect 435 706 437 716
rect 470 706 472 716
rect 581 706 583 716
rect 616 706 618 716
rect 747 706 749 716
rect 782 706 784 716
rect -330 674 -328 684
rect -295 674 -293 684
rect -260 674 -258 684
rect -164 674 -162 684
rect -129 674 -127 684
rect -27 674 -25 684
rect 8 674 10 684
rect 43 674 45 684
rect 139 674 141 684
rect 174 674 176 684
rect 269 674 271 684
rect 304 674 306 684
rect 339 674 341 684
rect 435 674 437 684
rect 470 674 472 684
rect 581 674 583 684
rect 616 674 618 684
rect 651 674 653 684
rect 747 674 749 684
rect 782 674 784 684
rect -279 -671 -277 -661
rect -244 -671 -242 -661
rect -113 -671 -111 -661
rect -78 -671 -76 -661
rect 24 -671 26 -661
rect 59 -671 61 -661
rect 190 -671 192 -661
rect 225 -671 227 -661
rect 320 -671 322 -661
rect 355 -671 357 -661
rect 486 -671 488 -661
rect 521 -671 523 -661
rect 632 -671 634 -661
rect 667 -671 669 -661
rect 798 -671 800 -661
rect 833 -671 835 -661
rect -279 -817 -277 -807
rect -244 -817 -242 -807
rect -113 -817 -111 -807
rect -78 -817 -76 -807
rect 24 -817 26 -807
rect 59 -817 61 -807
rect 190 -817 192 -807
rect 225 -817 227 -807
rect 320 -817 322 -807
rect 355 -817 357 -807
rect 486 -817 488 -807
rect 521 -817 523 -807
rect 632 -817 634 -807
rect 667 -817 669 -807
rect 798 -817 800 -807
rect 833 -817 835 -807
rect -279 -849 -277 -839
rect -244 -849 -242 -839
rect -209 -849 -207 -839
rect -113 -849 -111 -839
rect -78 -849 -76 -839
rect 24 -849 26 -839
rect 59 -849 61 -839
rect 94 -849 96 -839
rect 190 -849 192 -839
rect 225 -849 227 -839
rect 320 -849 322 -839
rect 355 -849 357 -839
rect 390 -849 392 -839
rect 486 -849 488 -839
rect 521 -849 523 -839
rect 632 -849 634 -839
rect 667 -849 669 -839
rect 702 -849 704 -839
rect 798 -849 800 -839
rect 833 -849 835 -839
<< ndiffusion >>
rect -313 817 -312 822
rect -310 817 -309 822
rect -147 817 -146 822
rect -144 817 -143 822
rect -10 817 -9 822
rect -7 817 -6 822
rect 156 817 157 822
rect 159 817 160 822
rect 286 817 287 822
rect 289 817 290 822
rect 452 817 453 822
rect 455 817 456 822
rect 598 817 599 822
rect 601 817 602 822
rect 764 817 765 822
rect 767 817 768 822
rect -313 797 -312 802
rect -310 797 -309 802
rect -147 797 -146 802
rect -144 797 -143 802
rect -10 797 -9 802
rect -7 797 -6 802
rect 156 797 157 802
rect 159 797 160 802
rect 286 797 287 802
rect 289 797 290 802
rect 452 797 453 802
rect 455 797 456 802
rect 598 797 599 802
rect 601 797 602 802
rect 764 797 765 802
rect 767 797 768 802
rect -313 766 -312 771
rect -310 766 -309 771
rect -147 766 -146 771
rect -144 766 -143 771
rect -10 766 -9 771
rect -7 766 -6 771
rect 156 766 157 771
rect 159 766 160 771
rect 286 766 287 771
rect 289 766 290 771
rect 452 766 453 771
rect 455 766 456 771
rect 598 766 599 771
rect 601 766 602 771
rect 764 766 765 771
rect 767 766 768 771
rect -313 746 -312 751
rect -310 746 -309 751
rect -147 746 -146 751
rect -144 746 -143 751
rect -10 746 -9 751
rect -7 746 -6 751
rect 156 746 157 751
rect 159 746 160 751
rect 286 746 287 751
rect 289 746 290 751
rect 452 746 453 751
rect 455 746 456 751
rect 598 746 599 751
rect 601 746 602 751
rect 764 746 765 751
rect 767 746 768 751
rect -313 639 -312 644
rect -310 639 -309 644
rect -313 615 -312 620
rect -310 615 -309 620
rect -147 639 -146 644
rect -144 639 -143 644
rect -10 639 -9 644
rect -7 639 -6 644
rect -147 619 -146 624
rect -144 619 -143 624
rect -10 615 -9 620
rect -7 615 -6 620
rect 156 639 157 644
rect 159 639 160 644
rect 286 639 287 644
rect 289 639 290 644
rect 156 619 157 624
rect 159 619 160 624
rect 286 615 287 620
rect 289 615 290 620
rect 452 639 453 644
rect 455 639 456 644
rect 598 639 599 644
rect 601 639 602 644
rect 452 619 453 624
rect 455 619 456 624
rect 598 615 599 620
rect 601 615 602 620
rect 764 639 765 644
rect 767 639 768 644
rect 764 619 765 624
rect 767 619 768 624
rect -313 596 -312 601
rect -310 596 -309 601
rect -10 596 -9 601
rect -7 596 -6 601
rect 286 596 287 601
rect 289 596 290 601
rect 598 596 599 601
rect 601 596 602 601
rect -262 -706 -261 -701
rect -259 -706 -258 -701
rect -96 -706 -95 -701
rect -93 -706 -92 -701
rect 41 -706 42 -701
rect 44 -706 45 -701
rect 207 -706 208 -701
rect 210 -706 211 -701
rect 337 -706 338 -701
rect 340 -706 341 -701
rect 503 -706 504 -701
rect 506 -706 507 -701
rect 649 -706 650 -701
rect 652 -706 653 -701
rect 815 -706 816 -701
rect 818 -706 819 -701
rect -262 -726 -261 -721
rect -259 -726 -258 -721
rect -96 -726 -95 -721
rect -93 -726 -92 -721
rect 41 -726 42 -721
rect 44 -726 45 -721
rect 207 -726 208 -721
rect 210 -726 211 -721
rect 337 -726 338 -721
rect 340 -726 341 -721
rect 503 -726 504 -721
rect 506 -726 507 -721
rect 649 -726 650 -721
rect 652 -726 653 -721
rect 815 -726 816 -721
rect 818 -726 819 -721
rect -262 -757 -261 -752
rect -259 -757 -258 -752
rect -96 -757 -95 -752
rect -93 -757 -92 -752
rect 41 -757 42 -752
rect 44 -757 45 -752
rect 207 -757 208 -752
rect 210 -757 211 -752
rect 337 -757 338 -752
rect 340 -757 341 -752
rect 503 -757 504 -752
rect 506 -757 507 -752
rect 649 -757 650 -752
rect 652 -757 653 -752
rect 815 -757 816 -752
rect 818 -757 819 -752
rect -262 -777 -261 -772
rect -259 -777 -258 -772
rect -96 -777 -95 -772
rect -93 -777 -92 -772
rect 41 -777 42 -772
rect 44 -777 45 -772
rect 207 -777 208 -772
rect 210 -777 211 -772
rect 337 -777 338 -772
rect 340 -777 341 -772
rect 503 -777 504 -772
rect 506 -777 507 -772
rect 649 -777 650 -772
rect 652 -777 653 -772
rect 815 -777 816 -772
rect 818 -777 819 -772
rect -262 -884 -261 -879
rect -259 -884 -258 -879
rect -262 -908 -261 -903
rect -259 -908 -258 -903
rect -96 -884 -95 -879
rect -93 -884 -92 -879
rect 41 -884 42 -879
rect 44 -884 45 -879
rect -96 -904 -95 -899
rect -93 -904 -92 -899
rect 41 -908 42 -903
rect 44 -908 45 -903
rect 207 -884 208 -879
rect 210 -884 211 -879
rect 337 -884 338 -879
rect 340 -884 341 -879
rect 207 -904 208 -899
rect 210 -904 211 -899
rect 337 -908 338 -903
rect 340 -908 341 -903
rect 503 -884 504 -879
rect 506 -884 507 -879
rect 649 -884 650 -879
rect 652 -884 653 -879
rect 503 -904 504 -899
rect 506 -904 507 -899
rect 649 -908 650 -903
rect 652 -908 653 -903
rect 815 -884 816 -879
rect 818 -884 819 -879
rect 815 -904 816 -899
rect 818 -904 819 -899
rect -262 -927 -261 -922
rect -259 -927 -258 -922
rect 41 -927 42 -922
rect 44 -927 45 -922
rect 337 -927 338 -922
rect 340 -927 341 -922
rect 649 -927 650 -922
rect 652 -927 653 -922
<< pdiffusion >>
rect -331 852 -330 862
rect -328 852 -327 862
rect -296 852 -295 862
rect -293 852 -292 862
rect -165 852 -164 862
rect -162 852 -161 862
rect -130 852 -129 862
rect -127 852 -126 862
rect -28 852 -27 862
rect -25 852 -24 862
rect 7 852 8 862
rect 10 852 11 862
rect 138 852 139 862
rect 141 852 142 862
rect 173 852 174 862
rect 176 852 177 862
rect 268 852 269 862
rect 271 852 272 862
rect 303 852 304 862
rect 306 852 307 862
rect 434 852 435 862
rect 437 852 438 862
rect 469 852 470 862
rect 472 852 473 862
rect 580 852 581 862
rect 583 852 584 862
rect 615 852 616 862
rect 618 852 619 862
rect 746 852 747 862
rect 749 852 750 862
rect 781 852 782 862
rect 784 852 785 862
rect -331 706 -330 716
rect -328 706 -327 716
rect -296 706 -295 716
rect -293 706 -292 716
rect -165 706 -164 716
rect -162 706 -161 716
rect -130 706 -129 716
rect -127 706 -126 716
rect -28 706 -27 716
rect -25 706 -24 716
rect 7 706 8 716
rect 10 706 11 716
rect 138 706 139 716
rect 141 706 142 716
rect 173 706 174 716
rect 176 706 177 716
rect 268 706 269 716
rect 271 706 272 716
rect 303 706 304 716
rect 306 706 307 716
rect 434 706 435 716
rect 437 706 438 716
rect 469 706 470 716
rect 472 706 473 716
rect 580 706 581 716
rect 583 706 584 716
rect 615 706 616 716
rect 618 706 619 716
rect 746 706 747 716
rect 749 706 750 716
rect 781 706 782 716
rect 784 706 785 716
rect -331 674 -330 684
rect -328 674 -327 684
rect -296 674 -295 684
rect -293 674 -292 684
rect -261 674 -260 684
rect -258 674 -257 684
rect -165 674 -164 684
rect -162 674 -161 684
rect -130 674 -129 684
rect -127 674 -126 684
rect -28 674 -27 684
rect -25 674 -24 684
rect 7 674 8 684
rect 10 674 11 684
rect 42 674 43 684
rect 45 674 46 684
rect 138 674 139 684
rect 141 674 142 684
rect 173 674 174 684
rect 176 674 177 684
rect 268 674 269 684
rect 271 674 272 684
rect 303 674 304 684
rect 306 674 307 684
rect 338 674 339 684
rect 341 674 342 684
rect 434 674 435 684
rect 437 674 438 684
rect 469 674 470 684
rect 472 674 473 684
rect 580 674 581 684
rect 583 674 584 684
rect 615 674 616 684
rect 618 674 619 684
rect 650 674 651 684
rect 653 674 654 684
rect 746 674 747 684
rect 749 674 750 684
rect 781 674 782 684
rect 784 674 785 684
rect -280 -671 -279 -661
rect -277 -671 -276 -661
rect -245 -671 -244 -661
rect -242 -671 -241 -661
rect -114 -671 -113 -661
rect -111 -671 -110 -661
rect -79 -671 -78 -661
rect -76 -671 -75 -661
rect 23 -671 24 -661
rect 26 -671 27 -661
rect 58 -671 59 -661
rect 61 -671 62 -661
rect 189 -671 190 -661
rect 192 -671 193 -661
rect 224 -671 225 -661
rect 227 -671 228 -661
rect 319 -671 320 -661
rect 322 -671 323 -661
rect 354 -671 355 -661
rect 357 -671 358 -661
rect 485 -671 486 -661
rect 488 -671 489 -661
rect 520 -671 521 -661
rect 523 -671 524 -661
rect 631 -671 632 -661
rect 634 -671 635 -661
rect 666 -671 667 -661
rect 669 -671 670 -661
rect 797 -671 798 -661
rect 800 -671 801 -661
rect 832 -671 833 -661
rect 835 -671 836 -661
rect -280 -817 -279 -807
rect -277 -817 -276 -807
rect -245 -817 -244 -807
rect -242 -817 -241 -807
rect -114 -817 -113 -807
rect -111 -817 -110 -807
rect -79 -817 -78 -807
rect -76 -817 -75 -807
rect 23 -817 24 -807
rect 26 -817 27 -807
rect 58 -817 59 -807
rect 61 -817 62 -807
rect 189 -817 190 -807
rect 192 -817 193 -807
rect 224 -817 225 -807
rect 227 -817 228 -807
rect 319 -817 320 -807
rect 322 -817 323 -807
rect 354 -817 355 -807
rect 357 -817 358 -807
rect 485 -817 486 -807
rect 488 -817 489 -807
rect 520 -817 521 -807
rect 523 -817 524 -807
rect 631 -817 632 -807
rect 634 -817 635 -807
rect 666 -817 667 -807
rect 669 -817 670 -807
rect 797 -817 798 -807
rect 800 -817 801 -807
rect 832 -817 833 -807
rect 835 -817 836 -807
rect -280 -849 -279 -839
rect -277 -849 -276 -839
rect -245 -849 -244 -839
rect -242 -849 -241 -839
rect -210 -849 -209 -839
rect -207 -849 -206 -839
rect -114 -849 -113 -839
rect -111 -849 -110 -839
rect -79 -849 -78 -839
rect -76 -849 -75 -839
rect 23 -849 24 -839
rect 26 -849 27 -839
rect 58 -849 59 -839
rect 61 -849 62 -839
rect 93 -849 94 -839
rect 96 -849 97 -839
rect 189 -849 190 -839
rect 192 -849 193 -839
rect 224 -849 225 -839
rect 227 -849 228 -839
rect 319 -849 320 -839
rect 322 -849 323 -839
rect 354 -849 355 -839
rect 357 -849 358 -839
rect 389 -849 390 -839
rect 392 -849 393 -839
rect 485 -849 486 -839
rect 488 -849 489 -839
rect 520 -849 521 -839
rect 523 -849 524 -839
rect 631 -849 632 -839
rect 634 -849 635 -839
rect 666 -849 667 -839
rect 669 -849 670 -839
rect 701 -849 702 -839
rect 704 -849 705 -839
rect 797 -849 798 -839
rect 800 -849 801 -839
rect 832 -849 833 -839
rect 835 -849 836 -839
<< ndcontact >>
rect -317 817 -313 822
rect -309 817 -305 822
rect -151 817 -147 822
rect -143 817 -139 822
rect -14 817 -10 822
rect -6 817 -2 822
rect 152 817 156 822
rect 160 817 164 822
rect 282 817 286 822
rect 290 817 294 822
rect 448 817 452 822
rect 456 817 460 822
rect 594 817 598 822
rect 602 817 606 822
rect 760 817 764 822
rect 768 817 772 822
rect -317 797 -313 802
rect -309 797 -305 802
rect -151 797 -147 802
rect -143 797 -139 802
rect -14 797 -10 802
rect -6 797 -2 802
rect 152 797 156 802
rect 160 797 164 802
rect 282 797 286 802
rect 290 797 294 802
rect 448 797 452 802
rect 456 797 460 802
rect 594 797 598 802
rect 602 797 606 802
rect 760 797 764 802
rect 768 797 772 802
rect -317 766 -313 771
rect -309 766 -305 771
rect -151 766 -147 771
rect -143 766 -139 771
rect -14 766 -10 771
rect -6 766 -2 771
rect 152 766 156 771
rect 160 766 164 771
rect 282 766 286 771
rect 290 766 294 771
rect 448 766 452 771
rect 456 766 460 771
rect 594 766 598 771
rect 602 766 606 771
rect 760 766 764 771
rect 768 766 772 771
rect -317 746 -313 751
rect -309 746 -305 751
rect -151 746 -147 751
rect -143 746 -139 751
rect -14 746 -10 751
rect -6 746 -2 751
rect 152 746 156 751
rect 160 746 164 751
rect 282 746 286 751
rect 290 746 294 751
rect 448 746 452 751
rect 456 746 460 751
rect 594 746 598 751
rect 602 746 606 751
rect 760 746 764 751
rect 768 746 772 751
rect -317 639 -313 644
rect -309 639 -305 644
rect -317 615 -313 620
rect -309 615 -305 620
rect -151 639 -147 644
rect -143 639 -139 644
rect -14 639 -10 644
rect -6 639 -2 644
rect -151 619 -147 624
rect -143 619 -139 624
rect -14 615 -10 620
rect -6 615 -2 620
rect 152 639 156 644
rect 160 639 164 644
rect 282 639 286 644
rect 290 639 294 644
rect 152 619 156 624
rect 160 619 164 624
rect 282 615 286 620
rect 290 615 294 620
rect 448 639 452 644
rect 456 639 460 644
rect 594 639 598 644
rect 602 639 606 644
rect 448 619 452 624
rect 456 619 460 624
rect 594 615 598 620
rect 602 615 606 620
rect 760 639 764 644
rect 768 639 772 644
rect 760 619 764 624
rect 768 619 772 624
rect -317 596 -313 601
rect -309 596 -305 601
rect -14 596 -10 601
rect -6 596 -2 601
rect 282 596 286 601
rect 290 596 294 601
rect 594 596 598 601
rect 602 596 606 601
rect -266 -706 -262 -701
rect -258 -706 -254 -701
rect -100 -706 -96 -701
rect -92 -706 -88 -701
rect 37 -706 41 -701
rect 45 -706 49 -701
rect 203 -706 207 -701
rect 211 -706 215 -701
rect 333 -706 337 -701
rect 341 -706 345 -701
rect 499 -706 503 -701
rect 507 -706 511 -701
rect 645 -706 649 -701
rect 653 -706 657 -701
rect 811 -706 815 -701
rect 819 -706 823 -701
rect -266 -726 -262 -721
rect -258 -726 -254 -721
rect -100 -726 -96 -721
rect -92 -726 -88 -721
rect 37 -726 41 -721
rect 45 -726 49 -721
rect 203 -726 207 -721
rect 211 -726 215 -721
rect 333 -726 337 -721
rect 341 -726 345 -721
rect 499 -726 503 -721
rect 507 -726 511 -721
rect 645 -726 649 -721
rect 653 -726 657 -721
rect 811 -726 815 -721
rect 819 -726 823 -721
rect -266 -757 -262 -752
rect -258 -757 -254 -752
rect -100 -757 -96 -752
rect -92 -757 -88 -752
rect 37 -757 41 -752
rect 45 -757 49 -752
rect 203 -757 207 -752
rect 211 -757 215 -752
rect 333 -757 337 -752
rect 341 -757 345 -752
rect 499 -757 503 -752
rect 507 -757 511 -752
rect 645 -757 649 -752
rect 653 -757 657 -752
rect 811 -757 815 -752
rect 819 -757 823 -752
rect -266 -777 -262 -772
rect -258 -777 -254 -772
rect -100 -777 -96 -772
rect -92 -777 -88 -772
rect 37 -777 41 -772
rect 45 -777 49 -772
rect 203 -777 207 -772
rect 211 -777 215 -772
rect 333 -777 337 -772
rect 341 -777 345 -772
rect 499 -777 503 -772
rect 507 -777 511 -772
rect 645 -777 649 -772
rect 653 -777 657 -772
rect 811 -777 815 -772
rect 819 -777 823 -772
rect -266 -884 -262 -879
rect -258 -884 -254 -879
rect -266 -908 -262 -903
rect -258 -908 -254 -903
rect -100 -884 -96 -879
rect -92 -884 -88 -879
rect 37 -884 41 -879
rect 45 -884 49 -879
rect -100 -904 -96 -899
rect -92 -904 -88 -899
rect 37 -908 41 -903
rect 45 -908 49 -903
rect 203 -884 207 -879
rect 211 -884 215 -879
rect 333 -884 337 -879
rect 341 -884 345 -879
rect 203 -904 207 -899
rect 211 -904 215 -899
rect 333 -908 337 -903
rect 341 -908 345 -903
rect 499 -884 503 -879
rect 507 -884 511 -879
rect 645 -884 649 -879
rect 653 -884 657 -879
rect 499 -904 503 -899
rect 507 -904 511 -899
rect 645 -908 649 -903
rect 653 -908 657 -903
rect 811 -884 815 -879
rect 819 -884 823 -879
rect 811 -904 815 -899
rect 819 -904 823 -899
rect -266 -927 -262 -922
rect -258 -927 -254 -922
rect 37 -927 41 -922
rect 45 -927 49 -922
rect 333 -927 337 -922
rect 341 -927 345 -922
rect 645 -927 649 -922
rect 653 -927 657 -922
<< pdcontact >>
rect -335 852 -331 862
rect -327 852 -323 862
rect -300 852 -296 862
rect -292 852 -288 862
rect -169 852 -165 862
rect -161 852 -157 862
rect -134 852 -130 862
rect -126 852 -122 862
rect -32 852 -28 862
rect -24 852 -20 862
rect 3 852 7 862
rect 11 852 15 862
rect 134 852 138 862
rect 142 852 146 862
rect 169 852 173 862
rect 177 852 181 862
rect 264 852 268 862
rect 272 852 276 862
rect 299 852 303 862
rect 307 852 311 862
rect 430 852 434 862
rect 438 852 442 862
rect 465 852 469 862
rect 473 852 477 862
rect 576 852 580 862
rect 584 852 588 862
rect 611 852 615 862
rect 619 852 623 862
rect 742 852 746 862
rect 750 852 754 862
rect 777 852 781 862
rect 785 852 789 862
rect -335 706 -331 716
rect -327 706 -323 716
rect -300 706 -296 716
rect -292 706 -288 716
rect -169 706 -165 716
rect -161 706 -157 716
rect -134 706 -130 716
rect -126 706 -122 716
rect -32 706 -28 716
rect -24 706 -20 716
rect 3 706 7 716
rect 11 706 15 716
rect 134 706 138 716
rect 142 706 146 716
rect 169 706 173 716
rect 177 706 181 716
rect 264 706 268 716
rect 272 706 276 716
rect 299 706 303 716
rect 307 706 311 716
rect 430 706 434 716
rect 438 706 442 716
rect 465 706 469 716
rect 473 706 477 716
rect 576 706 580 716
rect 584 706 588 716
rect 611 706 615 716
rect 619 706 623 716
rect 742 706 746 716
rect 750 706 754 716
rect 777 706 781 716
rect 785 706 789 716
rect -335 674 -331 684
rect -327 674 -323 684
rect -300 674 -296 684
rect -292 674 -288 684
rect -265 674 -261 684
rect -257 674 -253 684
rect -169 674 -165 684
rect -161 674 -157 684
rect -134 674 -130 684
rect -126 674 -122 684
rect -32 674 -28 684
rect -24 674 -20 684
rect 3 674 7 684
rect 11 674 15 684
rect 38 674 42 684
rect 46 674 50 684
rect 134 674 138 684
rect 142 674 146 684
rect 169 674 173 684
rect 177 674 181 684
rect 264 674 268 684
rect 272 674 276 684
rect 299 674 303 684
rect 307 674 311 684
rect 334 674 338 684
rect 342 674 346 684
rect 430 674 434 684
rect 438 674 442 684
rect 465 674 469 684
rect 473 674 477 684
rect 576 674 580 684
rect 584 674 588 684
rect 611 674 615 684
rect 619 674 623 684
rect 646 674 650 684
rect 654 674 658 684
rect 742 674 746 684
rect 750 674 754 684
rect 777 674 781 684
rect 785 674 789 684
rect -284 -671 -280 -661
rect -276 -671 -272 -661
rect -249 -671 -245 -661
rect -241 -671 -237 -661
rect -118 -671 -114 -661
rect -110 -671 -106 -661
rect -83 -671 -79 -661
rect -75 -671 -71 -661
rect 19 -671 23 -661
rect 27 -671 31 -661
rect 54 -671 58 -661
rect 62 -671 66 -661
rect 185 -671 189 -661
rect 193 -671 197 -661
rect 220 -671 224 -661
rect 228 -671 232 -661
rect 315 -671 319 -661
rect 323 -671 327 -661
rect 350 -671 354 -661
rect 358 -671 362 -661
rect 481 -671 485 -661
rect 489 -671 493 -661
rect 516 -671 520 -661
rect 524 -671 528 -661
rect 627 -671 631 -661
rect 635 -671 639 -661
rect 662 -671 666 -661
rect 670 -671 674 -661
rect 793 -671 797 -661
rect 801 -671 805 -661
rect 828 -671 832 -661
rect 836 -671 840 -661
rect -284 -817 -280 -807
rect -276 -817 -272 -807
rect -249 -817 -245 -807
rect -241 -817 -237 -807
rect -118 -817 -114 -807
rect -110 -817 -106 -807
rect -83 -817 -79 -807
rect -75 -817 -71 -807
rect 19 -817 23 -807
rect 27 -817 31 -807
rect 54 -817 58 -807
rect 62 -817 66 -807
rect 185 -817 189 -807
rect 193 -817 197 -807
rect 220 -817 224 -807
rect 228 -817 232 -807
rect 315 -817 319 -807
rect 323 -817 327 -807
rect 350 -817 354 -807
rect 358 -817 362 -807
rect 481 -817 485 -807
rect 489 -817 493 -807
rect 516 -817 520 -807
rect 524 -817 528 -807
rect 627 -817 631 -807
rect 635 -817 639 -807
rect 662 -817 666 -807
rect 670 -817 674 -807
rect 793 -817 797 -807
rect 801 -817 805 -807
rect 828 -817 832 -807
rect 836 -817 840 -807
rect -284 -849 -280 -839
rect -276 -849 -272 -839
rect -249 -849 -245 -839
rect -241 -849 -237 -839
rect -214 -849 -210 -839
rect -206 -849 -202 -839
rect -118 -849 -114 -839
rect -110 -849 -106 -839
rect -83 -849 -79 -839
rect -75 -849 -71 -839
rect 19 -849 23 -839
rect 27 -849 31 -839
rect 54 -849 58 -839
rect 62 -849 66 -839
rect 89 -849 93 -839
rect 97 -849 101 -839
rect 185 -849 189 -839
rect 193 -849 197 -839
rect 220 -849 224 -839
rect 228 -849 232 -839
rect 315 -849 319 -839
rect 323 -849 327 -839
rect 350 -849 354 -839
rect 358 -849 362 -839
rect 385 -849 389 -839
rect 393 -849 397 -839
rect 481 -849 485 -839
rect 489 -849 493 -839
rect 516 -849 520 -839
rect 524 -849 528 -839
rect 627 -849 631 -839
rect 635 -849 639 -839
rect 662 -849 666 -839
rect 670 -849 674 -839
rect 697 -849 701 -839
rect 705 -849 709 -839
rect 793 -849 797 -839
rect 801 -849 805 -839
rect 828 -849 832 -839
rect 836 -849 840 -839
<< polysilicon >>
rect -330 868 -284 870
rect -330 862 -328 868
rect -295 862 -293 865
rect -330 848 -328 852
rect -339 844 -328 848
rect -295 840 -293 852
rect -339 836 -293 840
rect -312 822 -310 836
rect -312 811 -310 817
rect -286 808 -284 868
rect -164 868 -118 870
rect -164 862 -162 868
rect -129 862 -127 865
rect -164 848 -162 852
rect -173 844 -162 848
rect -129 840 -127 852
rect -173 836 -127 840
rect -146 822 -144 836
rect -146 811 -144 817
rect -120 808 -118 868
rect -27 868 19 870
rect -27 862 -25 868
rect 8 862 10 865
rect -27 848 -25 852
rect -36 844 -25 848
rect 8 840 10 852
rect -36 836 10 840
rect -9 822 -7 836
rect -9 811 -7 817
rect 17 808 19 868
rect 139 868 185 870
rect 139 862 141 868
rect 174 862 176 865
rect 139 848 141 852
rect 130 844 141 848
rect 174 840 176 852
rect 130 836 176 840
rect 157 822 159 836
rect 157 811 159 817
rect 183 808 185 868
rect 269 868 315 870
rect 269 862 271 868
rect 304 862 306 865
rect 269 848 271 852
rect 260 844 271 848
rect 304 840 306 852
rect 260 836 306 840
rect 287 822 289 836
rect 287 811 289 817
rect 313 808 315 868
rect 435 868 481 870
rect 435 862 437 868
rect 470 862 472 865
rect 435 848 437 852
rect 426 844 437 848
rect 470 840 472 852
rect 426 836 472 840
rect 453 822 455 836
rect 453 811 455 817
rect 479 808 481 868
rect 581 868 627 870
rect 581 862 583 868
rect 616 862 618 865
rect 581 848 583 852
rect 572 844 583 848
rect 616 840 618 852
rect 572 836 618 840
rect 599 822 601 836
rect 599 811 601 817
rect 625 808 627 868
rect 747 868 793 870
rect 747 862 749 868
rect 782 862 784 865
rect 747 848 749 852
rect 738 844 749 848
rect 782 840 784 852
rect 738 836 784 840
rect 765 822 767 836
rect 765 811 767 817
rect 791 808 793 868
rect -312 806 -284 808
rect -146 806 -118 808
rect -9 806 19 808
rect 157 806 185 808
rect 287 806 315 808
rect 453 806 481 808
rect 599 806 627 808
rect 765 806 793 808
rect -312 802 -310 806
rect -146 802 -144 806
rect -9 802 -7 806
rect 157 802 159 806
rect 287 802 289 806
rect 453 802 455 806
rect 599 802 601 806
rect 765 802 767 806
rect -312 792 -310 797
rect -146 792 -144 797
rect -9 792 -7 797
rect 157 792 159 797
rect 287 792 289 797
rect 453 792 455 797
rect 599 792 601 797
rect 765 792 767 797
rect -312 771 -310 776
rect -146 771 -144 776
rect -9 771 -7 776
rect 157 771 159 776
rect 287 771 289 776
rect 453 771 455 776
rect 599 771 601 776
rect 765 771 767 776
rect -312 762 -310 766
rect -146 762 -144 766
rect -9 762 -7 766
rect 157 762 159 766
rect 287 762 289 766
rect 453 762 455 766
rect 599 762 601 766
rect 765 762 767 766
rect -312 760 -284 762
rect -146 760 -118 762
rect -9 760 19 762
rect 157 760 185 762
rect 287 760 315 762
rect 453 760 481 762
rect 599 760 627 762
rect 765 760 793 762
rect -312 751 -310 757
rect -312 732 -310 746
rect -339 728 -293 732
rect -339 720 -328 724
rect -330 716 -328 720
rect -295 716 -293 728
rect -330 700 -328 706
rect -295 703 -293 706
rect -286 700 -284 760
rect -146 751 -144 757
rect -146 732 -144 746
rect -173 728 -127 732
rect -173 720 -162 724
rect -164 716 -162 720
rect -129 716 -127 728
rect -330 698 -284 700
rect -164 700 -162 706
rect -129 703 -127 706
rect -120 700 -118 760
rect -9 751 -7 757
rect -9 732 -7 746
rect -36 728 10 732
rect -36 720 -25 724
rect -27 716 -25 720
rect 8 716 10 728
rect -164 698 -118 700
rect -27 700 -25 706
rect 8 703 10 706
rect 17 700 19 760
rect 157 751 159 757
rect 157 732 159 746
rect 130 728 176 732
rect 130 720 141 724
rect 139 716 141 720
rect 174 716 176 728
rect -27 698 19 700
rect 139 700 141 706
rect 174 703 176 706
rect 183 700 185 760
rect 287 751 289 757
rect 287 732 289 746
rect 260 728 306 732
rect 260 720 271 724
rect 269 716 271 720
rect 304 716 306 728
rect 139 698 185 700
rect 269 700 271 706
rect 304 703 306 706
rect 313 700 315 760
rect 453 751 455 757
rect 453 732 455 746
rect 426 728 472 732
rect 426 720 437 724
rect 435 716 437 720
rect 470 716 472 728
rect 269 698 315 700
rect 435 700 437 706
rect 470 703 472 706
rect 479 700 481 760
rect 599 751 601 757
rect 599 732 601 746
rect 572 728 618 732
rect 572 720 583 724
rect 581 716 583 720
rect 616 716 618 728
rect 435 698 481 700
rect 581 700 583 706
rect 616 703 618 706
rect 625 700 627 760
rect 765 751 767 757
rect 765 732 767 746
rect 738 728 784 732
rect 738 720 749 724
rect 747 716 749 720
rect 782 716 784 728
rect 581 698 627 700
rect 747 700 749 706
rect 782 703 784 706
rect 791 700 793 760
rect 747 698 793 700
rect -330 690 -284 692
rect -330 684 -328 690
rect -295 684 -293 687
rect -330 670 -328 674
rect -339 666 -328 670
rect -295 662 -293 674
rect -339 658 -293 662
rect -312 644 -310 658
rect -312 633 -310 639
rect -286 630 -284 690
rect -164 690 -118 692
rect -260 684 -258 687
rect -164 684 -162 690
rect -129 684 -127 687
rect -312 628 -284 630
rect -312 620 -310 628
rect -312 612 -310 615
rect -260 607 -258 674
rect -164 670 -162 674
rect -173 666 -162 670
rect -129 662 -127 674
rect -173 658 -127 662
rect -146 644 -144 658
rect -146 633 -144 639
rect -120 630 -118 690
rect -27 690 19 692
rect -27 684 -25 690
rect 8 684 10 687
rect -27 670 -25 674
rect -36 666 -25 670
rect 8 662 10 674
rect -36 658 10 662
rect -9 644 -7 658
rect -9 633 -7 639
rect 17 630 19 690
rect 139 690 185 692
rect 43 684 45 687
rect 139 684 141 690
rect 174 684 176 687
rect -146 628 -118 630
rect -9 628 19 630
rect -146 624 -144 628
rect -9 620 -7 628
rect -146 614 -144 619
rect -9 612 -7 615
rect 43 607 45 674
rect 139 670 141 674
rect 130 666 141 670
rect 174 662 176 674
rect 130 658 176 662
rect 157 644 159 658
rect 157 633 159 639
rect 183 630 185 690
rect 269 690 315 692
rect 269 684 271 690
rect 304 684 306 687
rect 269 670 271 674
rect 260 666 271 670
rect 304 662 306 674
rect 260 658 306 662
rect 287 644 289 658
rect 287 633 289 639
rect 313 630 315 690
rect 435 690 481 692
rect 339 684 341 687
rect 435 684 437 690
rect 470 684 472 687
rect 157 628 185 630
rect 287 628 315 630
rect 157 624 159 628
rect 287 620 289 628
rect 157 614 159 619
rect 287 612 289 615
rect 339 607 341 674
rect 435 670 437 674
rect 426 666 437 670
rect 470 662 472 674
rect 426 658 472 662
rect 453 644 455 658
rect 453 633 455 639
rect 479 630 481 690
rect 581 690 627 692
rect 581 684 583 690
rect 616 684 618 687
rect 581 670 583 674
rect 572 666 583 670
rect 616 662 618 674
rect 572 658 618 662
rect 599 644 601 658
rect 599 633 601 639
rect 625 630 627 690
rect 747 690 793 692
rect 651 684 653 687
rect 747 684 749 690
rect 782 684 784 687
rect 453 628 481 630
rect 599 628 627 630
rect 453 624 455 628
rect 599 620 601 628
rect 453 614 455 619
rect 599 612 601 615
rect 651 607 653 674
rect 747 670 749 674
rect 738 666 749 670
rect 782 662 784 674
rect 738 658 784 662
rect 765 644 767 658
rect 765 633 767 639
rect 791 630 793 690
rect 765 628 793 630
rect 765 624 767 628
rect 765 614 767 619
rect -312 605 -258 607
rect -9 605 45 607
rect 287 605 341 607
rect 599 605 653 607
rect -312 601 -310 605
rect -9 601 -7 605
rect 287 601 289 605
rect 599 601 601 605
rect -312 591 -310 596
rect -9 591 -7 596
rect 287 591 289 596
rect 599 591 601 596
rect -279 -655 -233 -653
rect -279 -661 -277 -655
rect -244 -661 -242 -658
rect -279 -675 -277 -671
rect -288 -679 -277 -675
rect -244 -683 -242 -671
rect -288 -687 -242 -683
rect -261 -701 -259 -687
rect -261 -712 -259 -706
rect -235 -715 -233 -655
rect -113 -655 -67 -653
rect -113 -661 -111 -655
rect -78 -661 -76 -658
rect -113 -675 -111 -671
rect -122 -679 -111 -675
rect -78 -683 -76 -671
rect -122 -687 -76 -683
rect -95 -701 -93 -687
rect -95 -712 -93 -706
rect -69 -715 -67 -655
rect 24 -655 70 -653
rect 24 -661 26 -655
rect 59 -661 61 -658
rect 24 -675 26 -671
rect 15 -679 26 -675
rect 59 -683 61 -671
rect 15 -687 61 -683
rect 42 -701 44 -687
rect 42 -712 44 -706
rect 68 -715 70 -655
rect 190 -655 236 -653
rect 190 -661 192 -655
rect 225 -661 227 -658
rect 190 -675 192 -671
rect 181 -679 192 -675
rect 225 -683 227 -671
rect 181 -687 227 -683
rect 208 -701 210 -687
rect 208 -712 210 -706
rect 234 -715 236 -655
rect 320 -655 366 -653
rect 320 -661 322 -655
rect 355 -661 357 -658
rect 320 -675 322 -671
rect 311 -679 322 -675
rect 355 -683 357 -671
rect 311 -687 357 -683
rect 338 -701 340 -687
rect 338 -712 340 -706
rect 364 -715 366 -655
rect 486 -655 532 -653
rect 486 -661 488 -655
rect 521 -661 523 -658
rect 486 -675 488 -671
rect 477 -679 488 -675
rect 521 -683 523 -671
rect 477 -687 523 -683
rect 504 -701 506 -687
rect 504 -712 506 -706
rect 530 -715 532 -655
rect 632 -655 678 -653
rect 632 -661 634 -655
rect 667 -661 669 -658
rect 632 -675 634 -671
rect 623 -679 634 -675
rect 667 -683 669 -671
rect 623 -687 669 -683
rect 650 -701 652 -687
rect 650 -712 652 -706
rect 676 -715 678 -655
rect 798 -655 844 -653
rect 798 -661 800 -655
rect 833 -661 835 -658
rect 798 -675 800 -671
rect 789 -679 800 -675
rect 833 -683 835 -671
rect 789 -687 835 -683
rect 816 -701 818 -687
rect 816 -712 818 -706
rect 842 -715 844 -655
rect -261 -717 -233 -715
rect -95 -717 -67 -715
rect 42 -717 70 -715
rect 208 -717 236 -715
rect 338 -717 366 -715
rect 504 -717 532 -715
rect 650 -717 678 -715
rect 816 -717 844 -715
rect -261 -721 -259 -717
rect -95 -721 -93 -717
rect 42 -721 44 -717
rect 208 -721 210 -717
rect 338 -721 340 -717
rect 504 -721 506 -717
rect 650 -721 652 -717
rect 816 -721 818 -717
rect -261 -731 -259 -726
rect -95 -731 -93 -726
rect 42 -731 44 -726
rect 208 -731 210 -726
rect 338 -731 340 -726
rect 504 -731 506 -726
rect 650 -731 652 -726
rect 816 -731 818 -726
rect -261 -752 -259 -747
rect -95 -752 -93 -747
rect 42 -752 44 -747
rect 208 -752 210 -747
rect 338 -752 340 -747
rect 504 -752 506 -747
rect 650 -752 652 -747
rect 816 -752 818 -747
rect -261 -761 -259 -757
rect -95 -761 -93 -757
rect 42 -761 44 -757
rect 208 -761 210 -757
rect 338 -761 340 -757
rect 504 -761 506 -757
rect 650 -761 652 -757
rect 816 -761 818 -757
rect -261 -763 -233 -761
rect -95 -763 -67 -761
rect 42 -763 70 -761
rect 208 -763 236 -761
rect 338 -763 366 -761
rect 504 -763 532 -761
rect 650 -763 678 -761
rect 816 -763 844 -761
rect -261 -772 -259 -766
rect -261 -791 -259 -777
rect -288 -795 -242 -791
rect -288 -803 -277 -799
rect -279 -807 -277 -803
rect -244 -807 -242 -795
rect -279 -823 -277 -817
rect -244 -820 -242 -817
rect -235 -823 -233 -763
rect -95 -772 -93 -766
rect -95 -791 -93 -777
rect -122 -795 -76 -791
rect -122 -803 -111 -799
rect -113 -807 -111 -803
rect -78 -807 -76 -795
rect -279 -825 -233 -823
rect -113 -823 -111 -817
rect -78 -820 -76 -817
rect -69 -823 -67 -763
rect 42 -772 44 -766
rect 42 -791 44 -777
rect 15 -795 61 -791
rect 15 -803 26 -799
rect 24 -807 26 -803
rect 59 -807 61 -795
rect -113 -825 -67 -823
rect 24 -823 26 -817
rect 59 -820 61 -817
rect 68 -823 70 -763
rect 208 -772 210 -766
rect 208 -791 210 -777
rect 181 -795 227 -791
rect 181 -803 192 -799
rect 190 -807 192 -803
rect 225 -807 227 -795
rect 24 -825 70 -823
rect 190 -823 192 -817
rect 225 -820 227 -817
rect 234 -823 236 -763
rect 338 -772 340 -766
rect 338 -791 340 -777
rect 311 -795 357 -791
rect 311 -803 322 -799
rect 320 -807 322 -803
rect 355 -807 357 -795
rect 190 -825 236 -823
rect 320 -823 322 -817
rect 355 -820 357 -817
rect 364 -823 366 -763
rect 504 -772 506 -766
rect 504 -791 506 -777
rect 477 -795 523 -791
rect 477 -803 488 -799
rect 486 -807 488 -803
rect 521 -807 523 -795
rect 320 -825 366 -823
rect 486 -823 488 -817
rect 521 -820 523 -817
rect 530 -823 532 -763
rect 650 -772 652 -766
rect 650 -791 652 -777
rect 623 -795 669 -791
rect 623 -803 634 -799
rect 632 -807 634 -803
rect 667 -807 669 -795
rect 486 -825 532 -823
rect 632 -823 634 -817
rect 667 -820 669 -817
rect 676 -823 678 -763
rect 816 -772 818 -766
rect 816 -791 818 -777
rect 789 -795 835 -791
rect 789 -803 800 -799
rect 798 -807 800 -803
rect 833 -807 835 -795
rect 632 -825 678 -823
rect 798 -823 800 -817
rect 833 -820 835 -817
rect 842 -823 844 -763
rect 798 -825 844 -823
rect -279 -833 -233 -831
rect -279 -839 -277 -833
rect -244 -839 -242 -836
rect -279 -853 -277 -849
rect -288 -857 -277 -853
rect -244 -861 -242 -849
rect -288 -865 -242 -861
rect -261 -879 -259 -865
rect -261 -890 -259 -884
rect -235 -893 -233 -833
rect -113 -833 -67 -831
rect -209 -839 -207 -836
rect -113 -839 -111 -833
rect -78 -839 -76 -836
rect -261 -895 -233 -893
rect -261 -903 -259 -895
rect -261 -911 -259 -908
rect -209 -916 -207 -849
rect -113 -853 -111 -849
rect -122 -857 -111 -853
rect -78 -861 -76 -849
rect -122 -865 -76 -861
rect -95 -879 -93 -865
rect -95 -890 -93 -884
rect -69 -893 -67 -833
rect 24 -833 70 -831
rect 24 -839 26 -833
rect 59 -839 61 -836
rect 24 -853 26 -849
rect 15 -857 26 -853
rect 59 -861 61 -849
rect 15 -865 61 -861
rect 42 -879 44 -865
rect 42 -890 44 -884
rect 68 -893 70 -833
rect 190 -833 236 -831
rect 94 -839 96 -836
rect 190 -839 192 -833
rect 225 -839 227 -836
rect -95 -895 -67 -893
rect 42 -895 70 -893
rect -95 -899 -93 -895
rect 42 -903 44 -895
rect -95 -909 -93 -904
rect 42 -911 44 -908
rect 94 -916 96 -849
rect 190 -853 192 -849
rect 181 -857 192 -853
rect 225 -861 227 -849
rect 181 -865 227 -861
rect 208 -879 210 -865
rect 208 -890 210 -884
rect 234 -893 236 -833
rect 320 -833 366 -831
rect 320 -839 322 -833
rect 355 -839 357 -836
rect 320 -853 322 -849
rect 311 -857 322 -853
rect 355 -861 357 -849
rect 311 -865 357 -861
rect 338 -879 340 -865
rect 338 -890 340 -884
rect 364 -893 366 -833
rect 486 -833 532 -831
rect 390 -839 392 -836
rect 486 -839 488 -833
rect 521 -839 523 -836
rect 208 -895 236 -893
rect 338 -895 366 -893
rect 208 -899 210 -895
rect 338 -903 340 -895
rect 208 -909 210 -904
rect 338 -911 340 -908
rect 390 -916 392 -849
rect 486 -853 488 -849
rect 477 -857 488 -853
rect 521 -861 523 -849
rect 477 -865 523 -861
rect 504 -879 506 -865
rect 504 -890 506 -884
rect 530 -893 532 -833
rect 632 -833 678 -831
rect 632 -839 634 -833
rect 667 -839 669 -836
rect 632 -853 634 -849
rect 623 -857 634 -853
rect 667 -861 669 -849
rect 623 -865 669 -861
rect 650 -879 652 -865
rect 650 -890 652 -884
rect 676 -893 678 -833
rect 798 -833 844 -831
rect 702 -839 704 -836
rect 798 -839 800 -833
rect 833 -839 835 -836
rect 504 -895 532 -893
rect 650 -895 678 -893
rect 504 -899 506 -895
rect 650 -903 652 -895
rect 504 -909 506 -904
rect 650 -911 652 -908
rect 702 -916 704 -849
rect 798 -853 800 -849
rect 789 -857 800 -853
rect 833 -861 835 -849
rect 789 -865 835 -861
rect 816 -879 818 -865
rect 816 -890 818 -884
rect 842 -893 844 -833
rect 816 -895 844 -893
rect 816 -899 818 -895
rect 816 -909 818 -904
rect -261 -918 -207 -916
rect 42 -918 96 -916
rect 338 -918 392 -916
rect 650 -918 704 -916
rect -261 -922 -259 -918
rect 42 -922 44 -918
rect 338 -922 340 -918
rect 650 -922 652 -918
rect -261 -932 -259 -927
rect 42 -932 44 -927
rect 338 -932 340 -927
rect 650 -932 652 -927
<< polycontact >>
rect -343 844 -339 848
rect -343 836 -339 840
rect -177 844 -173 848
rect -177 836 -173 840
rect -40 844 -36 848
rect -40 836 -36 840
rect 126 844 130 848
rect 126 836 130 840
rect 256 844 260 848
rect 256 836 260 840
rect 422 844 426 848
rect 422 836 426 840
rect 568 844 572 848
rect 568 836 572 840
rect 734 844 738 848
rect 734 836 738 840
rect -343 728 -339 732
rect -343 720 -339 724
rect -177 728 -173 732
rect -177 720 -173 724
rect -40 728 -36 732
rect -40 720 -36 724
rect 126 728 130 732
rect 126 720 130 724
rect 256 728 260 732
rect 256 720 260 724
rect 422 728 426 732
rect 422 720 426 724
rect 568 728 572 732
rect 568 720 572 724
rect 734 728 738 732
rect 734 720 738 724
rect -343 666 -339 670
rect -343 658 -339 662
rect -177 666 -173 670
rect -258 656 -254 660
rect -177 658 -173 662
rect -40 666 -36 670
rect -40 658 -36 662
rect 126 666 130 670
rect 45 656 49 660
rect 126 658 130 662
rect 256 666 260 670
rect 256 658 260 662
rect 422 666 426 670
rect 341 656 345 660
rect 422 658 426 662
rect 568 666 572 670
rect 568 658 572 662
rect 734 666 738 670
rect 653 656 657 660
rect 734 658 738 662
rect -292 -679 -288 -675
rect -292 -687 -288 -683
rect -126 -679 -122 -675
rect -126 -687 -122 -683
rect 11 -679 15 -675
rect 11 -687 15 -683
rect 177 -679 181 -675
rect 177 -687 181 -683
rect 307 -679 311 -675
rect 307 -687 311 -683
rect 473 -679 477 -675
rect 473 -687 477 -683
rect 619 -679 623 -675
rect 619 -687 623 -683
rect 785 -679 789 -675
rect 785 -687 789 -683
rect -292 -795 -288 -791
rect -292 -803 -288 -799
rect -126 -795 -122 -791
rect -126 -803 -122 -799
rect 11 -795 15 -791
rect 11 -803 15 -799
rect 177 -795 181 -791
rect 177 -803 181 -799
rect 307 -795 311 -791
rect 307 -803 311 -799
rect 473 -795 477 -791
rect 473 -803 477 -799
rect 619 -795 623 -791
rect 619 -803 623 -799
rect 785 -795 789 -791
rect 785 -803 789 -799
rect -292 -857 -288 -853
rect -292 -865 -288 -861
rect -126 -857 -122 -853
rect -207 -867 -203 -863
rect -126 -865 -122 -861
rect 11 -857 15 -853
rect 11 -865 15 -861
rect 177 -857 181 -853
rect 96 -867 100 -863
rect 177 -865 181 -861
rect 307 -857 311 -853
rect 307 -865 311 -861
rect 473 -857 477 -853
rect 392 -867 396 -863
rect 473 -865 477 -861
rect 619 -857 623 -853
rect 619 -865 623 -861
rect 785 -857 789 -853
rect 704 -867 708 -863
rect 785 -865 789 -861
<< metal1 >>
rect -341 870 795 873
rect -335 862 -331 870
rect -300 862 -296 870
rect -169 862 -165 870
rect -134 862 -130 870
rect -350 844 -348 849
rect -350 840 -343 841
rect -350 836 -348 840
rect -327 834 -323 852
rect -292 836 -288 852
rect -184 848 -177 849
rect -269 847 -177 848
rect -270 844 -177 847
rect -292 834 -282 836
rect -327 831 -282 834
rect -309 822 -305 831
rect -317 811 -313 817
rect -270 815 -265 844
rect -179 836 -177 841
rect -161 834 -157 852
rect -126 836 -122 852
rect -116 836 -111 841
rect -126 834 -116 836
rect -161 831 -116 834
rect -143 822 -139 831
rect -317 808 -305 811
rect -151 811 -147 817
rect -151 808 -139 811
rect -309 802 -305 808
rect -143 802 -139 808
rect -317 787 -313 797
rect -151 787 -147 797
rect -341 784 -263 787
rect -175 785 -116 787
rect -175 784 -123 785
rect -341 781 -123 784
rect -317 771 -313 781
rect -290 768 -277 773
rect -309 760 -305 766
rect -317 757 -305 760
rect -317 751 -313 757
rect -309 737 -305 746
rect -282 737 -277 768
rect -151 771 -147 781
rect -143 760 -139 766
rect -151 757 -139 760
rect -151 751 -147 757
rect -143 737 -139 746
rect -327 734 -282 737
rect -345 727 -343 732
rect -350 719 -343 724
rect -350 680 -346 719
rect -327 716 -323 734
rect -292 732 -282 734
rect -161 734 -116 737
rect -292 716 -288 732
rect -179 728 -177 732
rect -184 727 -177 728
rect -179 719 -177 724
rect -161 716 -157 734
rect -126 732 -116 734
rect -126 716 -122 732
rect -116 727 -111 732
rect -335 698 -331 706
rect -300 698 -296 706
rect -341 695 -282 698
rect -169 698 -165 706
rect -134 698 -130 706
rect -175 695 -116 698
rect -341 692 -116 695
rect -359 674 -346 680
rect -335 684 -331 692
rect -300 684 -296 692
rect -265 684 -261 692
rect -169 684 -165 692
rect -134 684 -130 692
rect -359 568 -356 674
rect -350 671 -346 674
rect -350 666 -343 671
rect -345 658 -343 663
rect -327 656 -323 674
rect -292 658 -288 674
rect -257 671 -253 674
rect -257 669 -235 671
rect -275 666 -235 669
rect -201 666 -184 671
rect -179 666 -177 671
rect -275 658 -271 666
rect -201 661 -196 666
rect -292 656 -271 658
rect -258 660 -247 661
rect -254 656 -247 660
rect -242 656 -196 661
rect -184 658 -177 663
rect -327 653 -271 656
rect -309 644 -305 653
rect -184 639 -179 658
rect -161 656 -157 674
rect -126 658 -122 674
rect -126 656 -116 658
rect -161 653 -116 656
rect -143 644 -139 653
rect -317 633 -313 639
rect -317 630 -305 633
rect -184 630 -179 634
rect -151 633 -147 639
rect -151 630 -139 633
rect -309 620 -305 630
rect -143 624 -139 630
rect -317 611 -313 615
rect -317 608 -305 611
rect -151 609 -147 619
rect -309 601 -305 608
rect -282 606 -116 609
rect -317 586 -313 596
rect -282 586 -279 606
rect -341 583 -279 586
rect -359 563 -101 568
rect -359 363 -356 563
rect -90 557 -87 870
rect -32 862 -28 870
rect 3 862 7 870
rect 134 862 138 870
rect 169 862 173 870
rect 264 862 268 870
rect 299 862 303 870
rect 430 862 434 870
rect 465 862 469 870
rect 576 862 580 870
rect 611 862 615 870
rect 742 862 746 870
rect 777 862 781 870
rect -47 844 -45 849
rect -47 840 -40 841
rect -47 836 -45 840
rect -24 834 -20 852
rect 11 836 15 852
rect 119 848 126 849
rect 34 847 126 848
rect 33 844 126 847
rect 11 834 21 836
rect -24 831 21 834
rect -6 822 -2 831
rect -14 811 -10 817
rect 33 815 38 844
rect 124 836 126 841
rect 142 834 146 852
rect 177 836 181 852
rect 249 844 251 849
rect 187 836 192 841
rect 249 840 256 841
rect 249 836 251 840
rect 177 834 187 836
rect 142 831 187 834
rect 272 834 276 852
rect 307 836 311 852
rect 415 848 422 849
rect 330 847 422 848
rect 329 844 422 847
rect 307 834 317 836
rect 272 831 317 834
rect 160 822 164 831
rect 290 822 294 831
rect -14 808 -2 811
rect 152 811 156 817
rect 282 811 286 817
rect 329 815 334 844
rect 420 836 422 841
rect 438 834 442 852
rect 473 836 477 852
rect 561 844 563 849
rect 483 836 488 841
rect 561 840 568 841
rect 561 836 563 840
rect 473 834 483 836
rect 438 831 483 834
rect 584 834 588 852
rect 619 836 623 852
rect 727 848 734 849
rect 642 847 734 848
rect 641 844 734 847
rect 619 834 629 836
rect 584 831 629 834
rect 456 822 460 831
rect 602 822 606 831
rect 152 808 164 811
rect 282 808 294 811
rect 448 811 452 817
rect 594 811 598 817
rect 641 815 646 844
rect 732 836 734 841
rect 750 834 754 852
rect 785 836 789 852
rect 795 836 800 841
rect 785 834 795 836
rect 750 831 795 834
rect 768 822 772 831
rect 448 808 460 811
rect 594 808 606 811
rect 760 811 764 817
rect 760 808 772 811
rect -6 802 -2 808
rect 160 802 164 808
rect 290 802 294 808
rect 456 802 460 808
rect 602 802 606 808
rect 768 802 772 808
rect -14 787 -10 797
rect 152 787 156 797
rect 282 787 286 797
rect 448 787 452 797
rect 594 787 598 797
rect 760 787 764 797
rect -38 786 40 787
rect -39 784 40 786
rect 128 784 336 787
rect 424 786 483 787
rect 570 786 648 787
rect 424 784 648 786
rect 736 784 795 787
rect -32 781 795 784
rect -32 778 -31 781
rect -14 771 -10 781
rect 13 768 26 773
rect -6 760 -2 766
rect -14 757 -2 760
rect -14 751 -10 757
rect -6 737 -2 746
rect 21 737 26 768
rect 152 771 156 781
rect 282 771 286 781
rect 309 768 322 773
rect 160 760 164 766
rect 290 760 294 766
rect 152 757 164 760
rect 282 757 294 760
rect 152 751 156 757
rect 282 751 286 757
rect 160 737 164 746
rect 290 737 294 746
rect 317 737 322 768
rect 448 771 452 781
rect 594 771 598 781
rect 621 768 634 773
rect 456 760 460 766
rect 602 760 606 766
rect 448 757 460 760
rect 594 757 606 760
rect 448 751 452 757
rect 594 751 598 757
rect 456 737 460 746
rect 602 737 606 746
rect 629 737 634 768
rect 760 771 764 781
rect 768 760 772 766
rect 760 757 772 760
rect 760 751 764 757
rect 768 737 772 746
rect -24 734 21 737
rect -42 727 -40 732
rect -47 719 -40 724
rect -47 676 -43 719
rect -24 716 -20 734
rect 11 732 21 734
rect 142 734 187 737
rect 11 716 15 732
rect 124 728 126 732
rect 119 727 126 728
rect 124 719 126 724
rect 142 716 146 734
rect 177 732 187 734
rect 272 734 317 737
rect 177 716 181 732
rect 187 727 192 732
rect 254 727 256 732
rect 249 719 256 724
rect -32 698 -28 706
rect 3 698 7 706
rect -38 695 21 698
rect 134 698 138 706
rect 169 698 173 706
rect 128 695 187 698
rect -38 692 187 695
rect -64 672 -43 676
rect -32 684 -28 692
rect 3 684 7 692
rect 38 684 42 692
rect 134 684 138 692
rect 169 684 173 692
rect 249 684 253 719
rect 272 716 276 734
rect 307 732 317 734
rect 438 734 483 737
rect 307 716 311 732
rect 420 728 422 732
rect 415 727 422 728
rect 420 719 422 724
rect 438 716 442 734
rect 473 732 483 734
rect 584 734 629 737
rect 473 716 477 732
rect 483 727 488 732
rect 566 727 568 732
rect 561 719 568 724
rect 264 698 268 706
rect 299 698 303 706
rect 258 695 317 698
rect 430 698 434 706
rect 465 698 469 706
rect 424 695 483 698
rect 258 692 483 695
rect -64 568 -60 672
rect -47 671 -43 672
rect -47 667 -40 671
rect -42 666 -40 667
rect -42 658 -40 663
rect -24 656 -20 674
rect 11 658 15 674
rect 46 671 50 674
rect 46 669 68 671
rect 28 666 68 669
rect 102 666 119 671
rect 124 666 126 671
rect 28 658 32 666
rect 102 661 107 666
rect 11 656 32 658
rect 45 660 56 661
rect 49 656 56 660
rect 61 656 107 661
rect 119 658 126 663
rect -24 653 32 656
rect -6 644 -2 653
rect 119 639 124 658
rect 142 656 146 674
rect 177 658 181 674
rect 239 678 253 684
rect 177 656 187 658
rect 142 653 187 656
rect 160 644 164 653
rect -14 633 -10 639
rect -14 630 -2 633
rect 119 630 124 634
rect 152 633 156 639
rect 152 630 164 633
rect -6 620 -2 630
rect 160 624 164 630
rect -14 611 -10 615
rect -14 608 -2 611
rect 152 609 156 619
rect -6 601 -2 608
rect 21 606 199 609
rect -14 586 -10 596
rect 21 586 24 606
rect -38 583 24 586
rect 239 568 243 678
rect 249 671 253 678
rect 264 684 268 692
rect 299 684 303 692
rect 334 684 338 692
rect 430 684 434 692
rect 465 684 469 692
rect 561 681 565 719
rect 584 716 588 734
rect 619 732 629 734
rect 750 734 795 737
rect 619 716 623 732
rect 732 728 734 732
rect 727 727 734 728
rect 732 719 734 724
rect 750 716 754 734
rect 785 732 795 734
rect 785 716 789 732
rect 795 727 800 732
rect 576 698 580 706
rect 611 698 615 706
rect 570 695 629 698
rect 742 698 746 706
rect 777 698 781 706
rect 736 695 795 698
rect 570 692 795 695
rect 249 666 256 671
rect 254 658 256 663
rect 272 656 276 674
rect 307 658 311 674
rect 342 671 346 674
rect 342 669 364 671
rect 324 666 364 669
rect 398 666 415 671
rect 420 666 422 671
rect 324 658 328 666
rect 398 661 403 666
rect 307 656 328 658
rect 341 660 352 661
rect 345 656 352 660
rect 357 656 403 661
rect 415 658 422 663
rect 272 653 328 656
rect 290 644 294 653
rect 415 639 420 658
rect 438 656 442 674
rect 473 658 477 674
rect 551 677 565 681
rect 473 656 483 658
rect 438 653 483 656
rect 456 644 460 653
rect 282 633 286 639
rect 282 630 294 633
rect 415 630 420 634
rect 448 633 452 639
rect 448 630 460 633
rect 290 620 294 630
rect 456 624 460 630
rect 282 611 286 615
rect 282 608 294 611
rect 448 609 452 619
rect 290 601 294 608
rect 317 606 487 609
rect 282 586 286 596
rect 317 586 320 606
rect 275 583 320 586
rect 551 568 555 677
rect 561 671 565 677
rect 576 684 580 692
rect 611 684 615 692
rect 646 684 650 692
rect 742 684 746 692
rect 777 684 781 692
rect 561 666 568 671
rect 566 658 568 663
rect 584 656 588 674
rect 619 658 623 674
rect 654 671 658 674
rect 654 669 676 671
rect 636 666 676 669
rect 710 666 727 671
rect 732 666 734 671
rect 636 658 640 666
rect 710 661 715 666
rect 619 656 640 658
rect 653 660 664 661
rect 657 656 664 660
rect 669 656 715 661
rect 727 658 734 663
rect 584 653 640 656
rect 602 644 606 653
rect 727 639 732 658
rect 750 656 754 674
rect 785 658 789 674
rect 785 656 795 658
rect 750 653 795 656
rect 768 644 772 653
rect 594 633 598 639
rect 594 630 606 633
rect 727 630 732 634
rect 760 633 764 639
rect 760 630 772 633
rect 602 620 606 630
rect 768 624 772 630
rect 594 611 598 615
rect 594 608 606 611
rect 760 609 764 619
rect 602 601 606 608
rect 629 606 795 609
rect 594 586 598 596
rect 629 586 632 606
rect 570 583 632 586
rect -76 563 555 568
rect 519 562 555 563
rect -118 554 -31 557
rect 184 554 271 557
rect 483 554 570 557
rect -117 469 -36 470
rect -117 465 -34 469
rect 187 465 268 469
rect 483 466 570 470
rect -117 464 -36 465
rect -120 377 -102 382
rect -116 376 -102 377
rect -184 314 -179 318
rect -124 168 -120 169
rect -107 168 -102 376
rect -56 358 -45 363
rect 238 362 251 367
rect 545 356 564 362
rect -47 179 -42 323
rect 119 314 124 318
rect 226 317 249 323
rect 125 223 129 291
rect 226 237 231 317
rect 415 314 420 318
rect 545 251 550 356
rect 727 314 732 318
rect 171 233 231 237
rect 42 208 47 222
rect 131 179 136 185
rect -47 174 136 179
rect 228 178 233 187
rect 176 173 233 178
rect 326 177 331 185
rect 291 172 331 177
rect 342 168 347 170
rect -124 165 12 168
rect -124 -34 -120 165
rect 361 71 364 72
rect 354 69 360 71
rect 136 -6 141 5
rect -100 -10 141 -6
rect 322 -52 327 -47
rect 322 -89 327 -57
rect 322 -93 334 -89
rect 378 -128 381 -58
rect -62 -215 -57 -179
rect -111 -262 50 -257
rect 303 -273 307 -224
rect 497 -273 598 -272
rect 390 -276 450 -273
rect 500 -275 598 -273
rect 558 -276 598 -275
rect 821 -307 826 -303
rect 500 -330 580 -326
rect 43 -335 48 -330
rect 2 -373 9 -370
rect 427 -373 487 -370
rect 500 -373 560 -370
rect 107 -505 117 -501
rect 215 -502 219 -501
rect 214 -505 219 -502
rect 317 -505 320 -501
rect 418 -502 419 -501
rect 417 -503 419 -502
rect 418 -504 419 -503
rect 417 -505 419 -504
rect 576 -505 580 -330
rect 821 -419 826 -415
rect 576 -511 590 -505
rect 219 -548 224 -545
rect 320 -548 325 -545
rect 419 -548 424 -545
rect -290 -653 459 -650
rect 464 -653 846 -650
rect -284 -661 -280 -653
rect -249 -661 -245 -653
rect -118 -661 -114 -653
rect -83 -661 -79 -653
rect 19 -661 23 -653
rect 54 -661 58 -653
rect 185 -661 189 -653
rect 220 -661 224 -653
rect 315 -661 319 -653
rect 350 -661 354 -653
rect 481 -661 485 -653
rect 516 -661 520 -653
rect 627 -661 631 -653
rect 662 -661 666 -653
rect 793 -661 797 -653
rect 828 -661 832 -653
rect -299 -679 -297 -674
rect -299 -683 -292 -682
rect -299 -687 -297 -683
rect -276 -689 -272 -671
rect -241 -687 -237 -671
rect -133 -675 -126 -674
rect -218 -676 -126 -675
rect -219 -679 -126 -676
rect -241 -689 -231 -687
rect -276 -692 -231 -689
rect -258 -701 -254 -692
rect -266 -712 -262 -706
rect -219 -708 -214 -679
rect -128 -687 -126 -682
rect -110 -689 -106 -671
rect -75 -687 -71 -671
rect 4 -679 6 -674
rect -65 -687 -60 -682
rect 4 -683 11 -682
rect 4 -687 6 -683
rect -75 -689 -65 -687
rect -110 -692 -65 -689
rect 27 -689 31 -671
rect 62 -687 66 -671
rect 170 -675 177 -674
rect 85 -676 177 -675
rect 84 -679 177 -676
rect 62 -689 72 -687
rect 27 -692 72 -689
rect -92 -701 -88 -692
rect 45 -701 49 -692
rect -266 -715 -254 -712
rect -100 -712 -96 -706
rect 37 -712 41 -706
rect 84 -708 89 -679
rect 175 -687 177 -682
rect 193 -689 197 -671
rect 228 -687 232 -671
rect 300 -679 302 -674
rect 238 -687 243 -682
rect 300 -683 307 -682
rect 300 -687 302 -683
rect 228 -689 238 -687
rect 193 -692 238 -689
rect 323 -689 327 -671
rect 358 -687 362 -671
rect 466 -675 473 -674
rect 381 -676 473 -675
rect 380 -679 473 -676
rect 358 -689 368 -687
rect 323 -692 368 -689
rect 211 -701 215 -692
rect 341 -701 345 -692
rect -100 -715 -88 -712
rect 37 -715 49 -712
rect 203 -712 207 -706
rect 333 -712 337 -706
rect 380 -708 385 -679
rect 471 -687 473 -682
rect 489 -689 493 -671
rect 524 -687 528 -671
rect 612 -679 614 -674
rect 534 -687 539 -682
rect 612 -683 619 -682
rect 612 -687 614 -683
rect 524 -689 534 -687
rect 489 -692 534 -689
rect 635 -689 639 -671
rect 670 -687 674 -671
rect 778 -675 785 -674
rect 693 -676 785 -675
rect 692 -679 785 -676
rect 670 -689 680 -687
rect 635 -692 680 -689
rect 507 -701 511 -692
rect 653 -701 657 -692
rect 203 -715 215 -712
rect 333 -715 345 -712
rect 499 -712 503 -706
rect 645 -712 649 -706
rect 692 -708 697 -679
rect 783 -687 785 -682
rect 801 -689 805 -671
rect 836 -687 840 -671
rect 846 -687 851 -682
rect 836 -689 846 -687
rect 801 -692 846 -689
rect 819 -701 823 -692
rect 499 -715 511 -712
rect 645 -715 657 -712
rect 811 -712 815 -706
rect 811 -715 823 -712
rect -258 -721 -254 -715
rect -92 -721 -88 -715
rect 45 -721 49 -715
rect 211 -721 215 -715
rect 341 -721 345 -715
rect 507 -721 511 -715
rect 653 -721 657 -715
rect 819 -721 823 -715
rect -266 -736 -262 -726
rect -100 -736 -96 -726
rect 37 -736 41 -726
rect 203 -736 207 -726
rect 333 -736 337 -726
rect 499 -736 503 -726
rect 645 -736 649 -726
rect 811 -736 815 -726
rect -290 -739 -212 -736
rect -124 -738 -65 -736
rect 13 -737 91 -736
rect -124 -739 -72 -738
rect -290 -742 -72 -739
rect -266 -752 -262 -742
rect -239 -755 -226 -750
rect -258 -763 -254 -757
rect -266 -766 -254 -763
rect -266 -772 -262 -766
rect -258 -786 -254 -777
rect -231 -786 -226 -755
rect -100 -752 -96 -742
rect 12 -739 91 -737
rect 179 -739 387 -736
rect 475 -737 534 -736
rect 621 -737 699 -736
rect 475 -739 699 -737
rect 787 -739 846 -736
rect 19 -742 846 -739
rect 19 -745 20 -742
rect 37 -752 41 -742
rect 64 -755 77 -750
rect -92 -763 -88 -757
rect 45 -763 49 -757
rect -100 -766 -88 -763
rect 37 -766 49 -763
rect -100 -772 -96 -766
rect 37 -772 41 -766
rect -92 -786 -88 -777
rect 45 -786 49 -777
rect 72 -786 77 -755
rect 203 -752 207 -742
rect 333 -752 337 -742
rect 360 -755 373 -750
rect 211 -763 215 -757
rect 341 -763 345 -757
rect 203 -766 215 -763
rect 333 -766 345 -763
rect 203 -772 207 -766
rect 333 -772 337 -766
rect 211 -786 215 -777
rect 341 -786 345 -777
rect 368 -786 373 -755
rect 499 -752 503 -742
rect 645 -752 649 -742
rect 672 -755 685 -750
rect 507 -763 511 -757
rect 653 -763 657 -757
rect 499 -766 511 -763
rect 645 -766 657 -763
rect 499 -772 503 -766
rect 645 -772 649 -766
rect 507 -786 511 -777
rect 653 -786 657 -777
rect 680 -786 685 -755
rect 811 -752 815 -742
rect 819 -763 823 -757
rect 811 -766 823 -763
rect 811 -772 815 -766
rect 819 -786 823 -777
rect -276 -789 -231 -786
rect -294 -796 -292 -791
rect -299 -804 -292 -799
rect -299 -843 -295 -804
rect -276 -807 -272 -789
rect -241 -791 -231 -789
rect -110 -789 -65 -786
rect -241 -807 -237 -791
rect -128 -795 -126 -791
rect -133 -796 -126 -795
rect -128 -804 -126 -799
rect -110 -807 -106 -789
rect -75 -791 -65 -789
rect 27 -789 72 -786
rect -75 -807 -71 -791
rect -65 -796 -60 -791
rect 9 -796 11 -791
rect 4 -804 11 -799
rect -284 -825 -280 -817
rect -249 -825 -245 -817
rect -290 -828 -231 -825
rect -118 -825 -114 -817
rect -83 -825 -79 -817
rect -124 -828 -65 -825
rect -290 -831 -65 -828
rect -303 -848 -295 -843
rect -308 -849 -295 -848
rect -284 -839 -280 -831
rect -249 -839 -245 -831
rect -214 -839 -210 -831
rect -118 -839 -114 -831
rect -83 -839 -79 -831
rect 4 -847 8 -804
rect 27 -807 31 -789
rect 62 -791 72 -789
rect 193 -789 238 -786
rect 62 -807 66 -791
rect 175 -795 177 -791
rect 170 -796 177 -795
rect 175 -804 177 -799
rect 193 -807 197 -789
rect 228 -791 238 -789
rect 323 -789 368 -786
rect 228 -807 232 -791
rect 238 -796 243 -791
rect 305 -796 307 -791
rect 300 -804 307 -799
rect 19 -825 23 -817
rect 54 -825 58 -817
rect 13 -828 72 -825
rect 185 -825 189 -817
rect 220 -825 224 -817
rect 179 -828 238 -825
rect 13 -831 238 -828
rect -308 -944 -305 -849
rect -299 -852 -295 -849
rect -299 -857 -292 -852
rect -294 -865 -292 -860
rect -276 -867 -272 -849
rect -241 -865 -237 -849
rect -206 -852 -202 -849
rect -206 -854 -184 -852
rect -224 -857 -184 -854
rect -150 -857 -133 -852
rect -128 -857 -126 -852
rect -224 -865 -220 -857
rect -150 -862 -145 -857
rect -241 -867 -220 -865
rect -207 -863 -196 -862
rect -203 -867 -196 -863
rect -191 -867 -145 -862
rect -133 -865 -126 -860
rect -276 -870 -220 -867
rect -258 -879 -254 -870
rect -133 -884 -128 -865
rect -110 -867 -106 -849
rect -75 -865 -71 -849
rect -13 -851 8 -847
rect 19 -839 23 -831
rect 54 -839 58 -831
rect 89 -839 93 -831
rect 185 -839 189 -831
rect 220 -839 224 -831
rect 300 -839 304 -804
rect 323 -807 327 -789
rect 358 -791 368 -789
rect 489 -789 534 -786
rect 358 -807 362 -791
rect 471 -795 473 -791
rect 466 -796 473 -795
rect 471 -804 473 -799
rect 489 -807 493 -789
rect 524 -791 534 -789
rect 635 -789 680 -786
rect 524 -807 528 -791
rect 534 -796 539 -791
rect 617 -796 619 -791
rect 612 -804 619 -799
rect 315 -825 319 -817
rect 350 -825 354 -817
rect 309 -828 368 -825
rect 481 -825 485 -817
rect 516 -825 520 -817
rect 475 -828 534 -825
rect 309 -831 534 -828
rect -75 -867 -65 -865
rect -110 -870 -65 -867
rect -92 -879 -88 -870
rect -266 -890 -262 -884
rect -100 -890 -96 -884
rect -266 -893 -254 -890
rect -100 -893 -88 -890
rect -258 -903 -254 -893
rect -92 -899 -88 -893
rect -266 -912 -262 -908
rect -266 -915 -254 -912
rect -100 -914 -96 -904
rect -258 -922 -254 -915
rect -231 -917 -65 -914
rect -266 -937 -262 -927
rect -231 -937 -228 -917
rect -290 -940 -228 -937
rect -13 -944 -9 -851
rect 4 -852 8 -851
rect 4 -857 11 -852
rect 9 -865 11 -860
rect 27 -867 31 -849
rect 62 -865 66 -849
rect 97 -852 101 -849
rect 97 -854 119 -852
rect 79 -857 119 -854
rect 153 -857 170 -852
rect 175 -857 177 -852
rect 79 -865 83 -857
rect 153 -862 158 -857
rect 62 -867 83 -865
rect 96 -863 107 -862
rect 100 -867 107 -863
rect 112 -867 158 -862
rect 170 -865 177 -860
rect 27 -870 83 -867
rect 45 -879 49 -870
rect 170 -884 175 -865
rect 193 -867 197 -849
rect 228 -865 232 -849
rect 290 -845 304 -839
rect 228 -867 238 -865
rect 193 -870 238 -867
rect 211 -879 215 -870
rect 37 -890 41 -884
rect 203 -890 207 -884
rect 37 -893 49 -890
rect 203 -893 215 -890
rect 45 -903 49 -893
rect 211 -899 215 -893
rect 37 -912 41 -908
rect 37 -915 49 -912
rect 203 -914 207 -904
rect 45 -922 49 -915
rect 72 -917 250 -914
rect 37 -937 41 -927
rect 72 -937 75 -917
rect 13 -940 75 -937
rect 290 -944 294 -845
rect 300 -852 304 -845
rect 315 -839 319 -831
rect 350 -839 354 -831
rect 385 -839 389 -831
rect 481 -839 485 -831
rect 516 -839 520 -831
rect 612 -842 616 -804
rect 635 -807 639 -789
rect 670 -791 680 -789
rect 801 -789 846 -786
rect 670 -807 674 -791
rect 783 -795 785 -791
rect 778 -796 785 -795
rect 783 -804 785 -799
rect 801 -807 805 -789
rect 836 -791 846 -789
rect 836 -807 840 -791
rect 846 -796 851 -791
rect 627 -825 631 -817
rect 662 -825 666 -817
rect 621 -828 680 -825
rect 793 -825 797 -817
rect 828 -825 832 -817
rect 787 -828 846 -825
rect 621 -831 846 -828
rect 300 -857 307 -852
rect 305 -865 307 -860
rect 323 -867 327 -849
rect 358 -865 362 -849
rect 393 -852 397 -849
rect 393 -854 415 -852
rect 375 -857 415 -854
rect 449 -857 466 -852
rect 471 -857 473 -852
rect 375 -865 379 -857
rect 449 -862 454 -857
rect 358 -867 379 -865
rect 392 -863 403 -862
rect 396 -867 403 -863
rect 408 -867 454 -862
rect 466 -865 473 -860
rect 323 -870 379 -867
rect 341 -879 345 -870
rect 466 -884 471 -865
rect 489 -867 493 -849
rect 524 -865 528 -849
rect 602 -846 616 -842
rect 524 -867 534 -865
rect 489 -870 534 -867
rect 507 -879 511 -870
rect 333 -890 337 -884
rect 499 -890 503 -884
rect 333 -893 345 -890
rect 499 -893 511 -890
rect 341 -903 345 -893
rect 507 -899 511 -893
rect 333 -912 337 -908
rect 333 -915 345 -912
rect 499 -914 503 -904
rect 341 -922 345 -915
rect 368 -917 538 -914
rect 333 -937 337 -927
rect 368 -937 371 -917
rect 326 -940 371 -937
rect -308 -947 557 -944
rect 602 -944 606 -846
rect 612 -852 616 -846
rect 627 -839 631 -831
rect 662 -839 666 -831
rect 697 -839 701 -831
rect 793 -839 797 -831
rect 828 -839 832 -831
rect 612 -857 619 -852
rect 617 -865 619 -860
rect 635 -867 639 -849
rect 670 -865 674 -849
rect 705 -852 709 -849
rect 705 -854 727 -852
rect 687 -857 727 -854
rect 761 -857 778 -852
rect 783 -857 785 -852
rect 687 -865 691 -857
rect 761 -862 766 -857
rect 670 -867 691 -865
rect 704 -863 715 -862
rect 708 -867 715 -863
rect 720 -867 766 -862
rect 778 -865 785 -860
rect 635 -870 691 -867
rect 653 -879 657 -870
rect 778 -884 783 -865
rect 801 -867 805 -849
rect 836 -865 840 -849
rect 836 -867 846 -865
rect 801 -870 846 -867
rect 819 -879 823 -870
rect 645 -890 649 -884
rect 811 -890 815 -884
rect 645 -893 657 -890
rect 811 -893 823 -890
rect 653 -903 657 -893
rect 819 -899 823 -893
rect 645 -912 649 -908
rect 645 -915 657 -912
rect 811 -914 815 -904
rect 653 -922 657 -915
rect 680 -917 846 -914
rect 645 -937 649 -927
rect 680 -937 683 -917
rect 621 -940 683 -937
rect 562 -947 606 -944
<< m2contact >>
rect -348 844 -343 849
rect -348 835 -343 840
rect -282 831 -277 836
rect -116 831 -111 836
rect -270 810 -265 815
rect -295 768 -290 773
rect -123 779 -116 785
rect -350 727 -345 732
rect -282 732 -277 737
rect -184 728 -179 733
rect -350 658 -345 663
rect -184 666 -179 671
rect -247 656 -242 661
rect -116 653 -111 658
rect -350 634 -345 639
rect -184 634 -179 639
rect -101 563 -96 568
rect -45 844 -40 849
rect -45 835 -40 840
rect 21 831 26 836
rect 251 844 256 849
rect 187 831 192 836
rect 251 835 256 840
rect 317 831 322 836
rect 33 810 38 815
rect 563 844 568 849
rect 483 831 488 836
rect 563 835 568 840
rect 629 831 634 836
rect 329 810 334 815
rect 795 831 800 836
rect 641 810 646 815
rect -39 778 -32 784
rect 8 768 13 773
rect 304 768 309 773
rect 616 768 621 773
rect -47 727 -42 732
rect 21 732 26 737
rect 119 728 124 733
rect 249 727 254 732
rect 317 732 322 737
rect 415 728 420 733
rect 561 727 566 732
rect -47 658 -42 663
rect 119 666 124 671
rect 56 656 61 661
rect 187 653 192 658
rect -47 634 -42 639
rect 119 634 124 639
rect 629 732 634 737
rect 727 728 732 733
rect 249 658 254 663
rect 415 666 420 671
rect 352 656 357 661
rect 483 653 488 658
rect 249 634 254 639
rect 415 634 420 639
rect 561 658 566 663
rect 727 666 732 671
rect 664 656 669 661
rect 795 653 800 658
rect 561 634 566 639
rect 727 634 732 639
rect -81 563 -76 568
rect -359 358 -350 363
rect -61 358 -56 363
rect 233 362 238 367
rect 42 222 47 227
rect 545 245 550 251
rect 137 211 142 216
rect 234 211 239 216
rect 286 172 291 177
rect 377 63 382 68
rect 233 0 238 5
rect 331 -1 336 4
rect -105 -11 -100 -6
rect 322 -47 327 -42
rect -105 -84 -100 -79
rect 377 -58 382 -53
rect 555 -56 560 -51
rect -163 -184 -158 -179
rect -62 -220 -57 -215
rect 446 -330 451 -325
rect 560 -373 565 -368
rect 596 -366 601 -361
rect 586 -457 591 -452
rect 459 -653 464 -648
rect -297 -679 -292 -674
rect -297 -688 -292 -683
rect -231 -692 -226 -687
rect 6 -679 11 -674
rect -65 -692 -60 -687
rect 6 -688 11 -683
rect 72 -692 77 -687
rect -219 -713 -214 -708
rect 302 -679 307 -674
rect 238 -692 243 -687
rect 302 -688 307 -683
rect 368 -692 373 -687
rect 84 -713 89 -708
rect 614 -679 619 -674
rect 534 -692 539 -687
rect 614 -688 619 -683
rect 680 -692 685 -687
rect 380 -713 385 -708
rect 846 -692 851 -687
rect 692 -713 697 -708
rect -244 -755 -239 -750
rect -72 -744 -65 -738
rect 12 -745 19 -739
rect 59 -755 64 -750
rect 355 -755 360 -750
rect 667 -755 672 -750
rect -299 -796 -294 -791
rect -231 -791 -226 -786
rect -133 -795 -128 -790
rect 4 -796 9 -791
rect -308 -848 -303 -843
rect 72 -791 77 -786
rect 170 -795 175 -790
rect 300 -796 305 -791
rect -299 -865 -294 -860
rect -133 -857 -128 -852
rect -196 -867 -191 -862
rect 368 -791 373 -786
rect 466 -795 471 -790
rect 612 -796 617 -791
rect -65 -870 -60 -865
rect -299 -889 -294 -884
rect -133 -889 -128 -884
rect 4 -865 9 -860
rect 170 -857 175 -852
rect 107 -867 112 -862
rect 238 -870 243 -865
rect 4 -889 9 -884
rect 170 -889 175 -884
rect 680 -791 685 -786
rect 778 -795 783 -790
rect 300 -865 305 -860
rect 466 -857 471 -852
rect 403 -867 408 -862
rect 534 -870 539 -865
rect 300 -889 305 -884
rect 466 -889 471 -884
rect 557 -947 562 -942
rect 612 -865 617 -860
rect 778 -857 783 -852
rect 715 -867 720 -862
rect 846 -870 851 -865
rect 612 -889 617 -884
rect 778 -889 783 -884
<< metal2 >>
rect -343 844 -226 849
rect -40 844 77 849
rect 256 844 373 849
rect 568 844 685 849
rect -348 791 -343 835
rect -348 788 -289 791
rect -295 773 -289 788
rect -282 763 -277 831
rect -350 759 -277 763
rect -350 732 -345 759
rect -270 737 -265 810
rect -277 732 -242 737
rect -350 652 -345 658
rect -247 661 -242 732
rect -230 698 -226 844
rect -116 792 -111 831
rect -184 789 -111 792
rect -45 791 -40 835
rect -184 733 -180 789
rect -45 788 14 791
rect -116 779 -39 783
rect 8 773 14 788
rect 21 763 26 831
rect -47 759 26 763
rect -47 732 -42 759
rect 33 737 38 810
rect 26 732 61 737
rect -230 693 -111 698
rect -194 652 -189 693
rect -116 658 -111 693
rect -350 649 -189 652
rect -47 652 -42 658
rect 56 661 61 732
rect 73 698 77 844
rect 187 792 192 831
rect 119 789 192 792
rect 251 791 256 835
rect 119 733 123 789
rect 251 788 310 791
rect 304 773 310 788
rect 317 763 322 831
rect 249 759 322 763
rect 249 732 254 759
rect 329 737 334 810
rect 322 732 357 737
rect 73 693 192 698
rect 109 652 114 693
rect 187 658 192 693
rect -47 649 114 652
rect 249 652 254 658
rect 352 661 357 732
rect 369 698 373 844
rect 483 792 488 831
rect 415 789 488 792
rect 563 791 568 835
rect 415 733 419 789
rect 563 788 622 791
rect 616 773 622 788
rect 629 763 634 831
rect 561 759 634 763
rect 561 732 566 759
rect 641 737 646 810
rect 634 732 669 737
rect 369 693 488 698
rect 405 652 410 693
rect 483 658 488 693
rect 249 649 410 652
rect 561 652 566 658
rect 664 661 669 732
rect 681 698 685 844
rect 795 792 800 831
rect 727 789 800 792
rect 727 733 731 789
rect 681 693 800 698
rect 717 652 722 693
rect 795 658 800 693
rect 561 649 722 652
rect -387 634 -350 639
rect -345 634 -184 639
rect -67 634 -47 639
rect -42 634 119 639
rect 221 634 249 639
rect 254 634 415 639
rect 533 634 561 639
rect 566 634 727 639
rect -96 563 -81 568
rect -421 363 -350 365
rect -421 358 -359 363
rect -421 251 -416 358
rect -350 260 -345 323
rect -61 251 -56 358
rect 233 251 238 362
rect -421 245 545 251
rect -421 -618 -416 245
rect 561 236 566 318
rect 286 231 566 236
rect -180 222 42 227
rect -180 -95 -174 222
rect 94 212 137 216
rect 94 -4 97 212
rect 189 211 234 216
rect 131 174 136 182
rect -105 -71 -100 -11
rect -111 -72 -100 -71
rect -105 -79 -100 -72
rect -36 -10 97 -4
rect -36 -93 -31 -10
rect 189 -11 193 211
rect 286 177 291 231
rect 176 -16 193 -11
rect 233 -25 238 0
rect 78 -28 238 -25
rect 322 -1 331 4
rect 78 -88 83 -28
rect 322 -42 327 -1
rect 377 -53 382 63
rect -163 -231 -158 -184
rect -57 -220 200 -216
rect -163 -236 105 -231
rect 100 -361 105 -236
rect 195 -361 200 -220
rect 555 -247 560 -56
rect 446 -251 560 -247
rect 446 -325 451 -251
rect 596 -368 601 -366
rect 565 -373 601 -368
rect 385 -434 463 -433
rect 385 -438 464 -434
rect 461 -602 464 -438
rect -421 -621 -302 -618
rect -308 -843 -303 -621
rect 459 -648 464 -602
rect 557 -457 586 -452
rect -292 -679 -175 -674
rect 11 -679 128 -674
rect 307 -679 424 -674
rect -297 -732 -292 -688
rect -297 -735 -238 -732
rect -244 -750 -238 -735
rect -231 -760 -226 -692
rect -299 -764 -226 -760
rect -299 -791 -294 -764
rect -219 -786 -214 -713
rect -226 -791 -191 -786
rect -299 -871 -294 -865
rect -196 -862 -191 -791
rect -179 -825 -175 -679
rect -65 -731 -60 -692
rect -133 -734 -60 -731
rect 6 -732 11 -688
rect -133 -790 -129 -734
rect 6 -735 65 -732
rect -65 -744 12 -740
rect -39 -745 -35 -744
rect 59 -750 65 -735
rect 72 -760 77 -692
rect 4 -764 77 -760
rect 4 -791 9 -764
rect 84 -786 89 -713
rect 77 -791 112 -786
rect -179 -830 -60 -825
rect -143 -871 -138 -830
rect -65 -865 -60 -830
rect -299 -874 -138 -871
rect 4 -871 9 -865
rect 107 -862 112 -791
rect 124 -825 128 -679
rect 238 -731 243 -692
rect 170 -734 243 -731
rect 302 -732 307 -688
rect 170 -790 174 -734
rect 302 -735 361 -732
rect 355 -750 361 -735
rect 368 -760 373 -692
rect 300 -764 373 -760
rect 300 -791 305 -764
rect 380 -786 385 -713
rect 373 -791 408 -786
rect 124 -830 243 -825
rect 160 -871 165 -830
rect 238 -865 243 -830
rect 4 -874 165 -871
rect 300 -871 305 -865
rect 403 -862 408 -791
rect 420 -825 424 -679
rect 534 -731 539 -692
rect 466 -734 539 -731
rect 466 -790 470 -734
rect 420 -830 539 -825
rect 456 -871 461 -830
rect 534 -865 539 -830
rect 300 -874 461 -871
rect -321 -889 -299 -884
rect -294 -889 -133 -884
rect -16 -889 4 -884
rect 9 -889 170 -884
rect 272 -889 300 -884
rect 305 -889 466 -884
rect 557 -942 561 -457
rect 619 -679 736 -674
rect 614 -732 619 -688
rect 614 -735 673 -732
rect 667 -750 673 -735
rect 680 -760 685 -692
rect 612 -764 685 -760
rect 612 -791 617 -764
rect 692 -786 697 -713
rect 685 -791 720 -786
rect 612 -871 617 -865
rect 715 -862 720 -791
rect 732 -825 736 -679
rect 846 -731 851 -692
rect 778 -734 851 -731
rect 778 -790 782 -734
rect 732 -830 851 -825
rect 768 -871 773 -830
rect 846 -865 851 -830
rect 612 -874 773 -871
rect 584 -889 612 -884
rect 617 -889 778 -884
<< m3contact >>
rect -392 634 -387 639
rect -72 634 -67 639
rect 216 634 221 639
rect 528 634 533 639
rect -350 255 -345 260
rect 36 147 41 152
rect -111 -71 -105 -66
rect 78 -146 83 -141
rect -326 -889 -321 -884
rect -21 -889 -16 -884
rect 267 -889 272 -884
rect 579 -889 584 -884
<< m123contact >>
rect -279 865 -274 870
rect 24 865 29 870
rect 320 865 325 870
rect 632 865 637 870
rect -247 776 -242 781
rect -279 695 -274 700
rect -184 836 -179 841
rect -116 732 -111 737
rect 56 776 61 781
rect -184 719 -179 724
rect 24 695 29 700
rect -235 666 -230 671
rect 119 836 124 841
rect 187 732 192 737
rect 352 776 357 781
rect 119 719 124 724
rect 320 695 325 700
rect 68 666 73 671
rect 415 836 420 841
rect 483 732 488 737
rect 664 776 669 781
rect 415 719 420 724
rect 632 695 637 700
rect 364 666 369 671
rect 727 836 732 841
rect 795 732 800 737
rect 727 719 732 724
rect 676 666 681 671
rect -247 609 -242 614
rect 56 609 61 614
rect 352 609 357 614
rect 664 609 669 614
rect 171 228 176 233
rect -1 106 4 111
rect 38 0 43 5
rect 171 173 176 178
rect 102 106 107 111
rect 332 211 337 216
rect 197 106 202 111
rect 295 106 300 111
rect 171 -16 176 -11
rect 322 -57 327 -52
rect 171 -92 176 -87
rect 505 -171 510 -166
rect -2 -180 3 -175
rect 227 -179 232 -174
rect -116 -262 -111 -257
rect 50 -262 55 -257
rect -2 -335 3 -330
rect 38 -335 43 -330
rect 142 -335 147 -330
rect 239 -335 244 -330
rect 293 -335 298 -330
rect 337 -335 342 -330
rect 117 -506 122 -501
rect 219 -506 224 -501
rect 320 -506 325 -501
rect 419 -506 424 -501
rect 256 -553 261 -548
rect -228 -658 -223 -653
rect 75 -658 80 -653
rect 371 -658 376 -653
rect -196 -747 -191 -742
rect -228 -828 -223 -823
rect -133 -687 -128 -682
rect -65 -791 -60 -786
rect 107 -747 112 -742
rect -133 -804 -128 -799
rect 75 -828 80 -823
rect -184 -857 -179 -852
rect 170 -687 175 -682
rect 238 -791 243 -786
rect 403 -747 408 -742
rect 170 -804 175 -799
rect 371 -828 376 -823
rect 119 -857 124 -852
rect 466 -687 471 -682
rect 534 -791 539 -786
rect 466 -804 471 -799
rect 415 -857 420 -852
rect -196 -914 -191 -909
rect 107 -914 112 -909
rect 403 -914 408 -909
rect 683 -658 688 -653
rect 715 -747 720 -742
rect 683 -828 688 -823
rect 778 -687 783 -682
rect 846 -791 851 -786
rect 778 -804 783 -799
rect 727 -857 732 -852
rect 715 -914 720 -909
<< metal3 >>
rect -279 836 -274 865
rect -282 831 -274 836
rect -279 700 -274 831
rect 24 836 29 865
rect -392 246 -388 634
rect -247 614 -242 776
rect -184 764 -179 836
rect 21 831 29 836
rect -184 761 -111 764
rect -116 737 -111 761
rect -235 719 -184 724
rect -179 719 -178 724
rect -235 671 -230 719
rect 24 700 29 831
rect 320 836 325 865
rect -345 255 -136 260
rect -392 242 -150 246
rect -154 111 -150 242
rect -141 152 -136 255
rect -72 246 -68 634
rect 56 614 61 776
rect 119 764 124 836
rect 317 831 325 836
rect 119 761 192 764
rect 187 737 192 761
rect 68 719 119 724
rect 124 719 125 724
rect 68 671 73 719
rect 320 700 325 831
rect 632 836 637 865
rect 216 247 220 634
rect 352 614 357 776
rect 415 764 420 836
rect 629 831 637 836
rect 415 761 488 764
rect 483 737 488 761
rect 364 719 415 724
rect 420 719 421 724
rect 364 671 369 719
rect 632 700 637 831
rect -72 242 107 246
rect -72 241 -68 242
rect -141 147 36 152
rect 102 111 107 242
rect 191 242 221 247
rect 171 178 176 228
rect -154 106 -1 111
rect 4 106 5 111
rect 191 111 196 242
rect 528 236 533 634
rect 664 614 669 776
rect 727 764 732 836
rect 727 761 800 764
rect 795 737 800 761
rect 676 719 727 724
rect 732 719 733 724
rect 676 671 681 719
rect 296 235 533 236
rect 295 231 533 235
rect 295 111 300 231
rect 528 230 533 231
rect 337 211 435 216
rect 191 106 197 111
rect -116 -257 -111 -66
rect 3 -180 4 -175
rect -2 -330 1 -180
rect 38 -330 42 0
rect 171 -87 176 -16
rect 327 -57 374 -52
rect 72 -146 78 -141
rect 72 -249 77 -146
rect 227 -240 232 -179
rect 369 -229 374 -57
rect 430 -166 435 211
rect 430 -171 505 -166
rect 337 -234 374 -229
rect 227 -244 298 -240
rect 72 -254 244 -249
rect 55 -262 147 -258
rect 142 -330 147 -262
rect 239 -330 244 -254
rect 293 -330 298 -244
rect 337 -330 342 -234
rect -247 -576 -242 -575
rect 117 -576 122 -506
rect -247 -577 122 -576
rect -326 -581 122 -577
rect -326 -582 -242 -581
rect -326 -884 -321 -582
rect 219 -591 224 -506
rect -21 -595 224 -591
rect -228 -687 -223 -658
rect -231 -692 -223 -687
rect -228 -823 -223 -692
rect -326 -890 -321 -889
rect -196 -909 -191 -747
rect -133 -759 -128 -687
rect -133 -762 -60 -759
rect -65 -786 -60 -762
rect -184 -804 -133 -799
rect -128 -804 -127 -799
rect -184 -852 -179 -804
rect -21 -884 -15 -595
rect 20 -596 224 -595
rect 256 -605 261 -553
rect 320 -554 325 -506
rect 107 -609 261 -605
rect 267 -560 325 -554
rect 419 -554 424 -506
rect 552 -554 584 -553
rect 419 -558 584 -554
rect 552 -559 584 -558
rect 267 -605 273 -560
rect 75 -687 80 -658
rect 72 -692 80 -687
rect 75 -823 80 -692
rect 107 -742 112 -609
rect 107 -909 112 -747
rect 170 -759 175 -687
rect 170 -762 243 -759
rect 238 -786 243 -762
rect 119 -804 170 -799
rect 175 -804 176 -799
rect 119 -852 124 -804
rect 267 -884 272 -605
rect 371 -687 376 -658
rect 368 -692 376 -687
rect 371 -823 376 -692
rect 403 -909 408 -747
rect 466 -759 471 -687
rect 466 -762 539 -759
rect 534 -786 539 -762
rect 415 -804 466 -799
rect 471 -804 472 -799
rect 415 -852 420 -804
rect 579 -884 584 -559
rect 683 -687 688 -658
rect 680 -692 688 -687
rect 683 -823 688 -692
rect 579 -890 584 -889
rect 715 -909 720 -747
rect 778 -759 783 -687
rect 778 -762 851 -759
rect 846 -786 851 -762
rect 727 -804 778 -799
rect 783 -804 784 -799
rect 727 -852 732 -804
use dff  dff_0
timestamp 1619465570
transform 1 0 -350 0 1 468
box 0 -201 239 89
use dff  dff_1
timestamp 1619465570
transform 1 0 -47 0 1 468
box 0 -201 239 89
use dff  dff_2
timestamp 1619465570
transform 1 0 249 0 1 468
box 0 -201 239 89
use dff  dff_3
timestamp 1619465570
transform 1 0 561 0 1 468
box 0 -201 239 89
use pg  pg_0
timestamp 1619529852
transform 1 0 9 0 1 68
box -9 -68 382 155
use cla  cla_0
timestamp 1619529852
transform 1 0 -171 0 1 -131
box -20 -95 741 100
use sum  sum_0
timestamp 1619527417
transform 1 0 7 0 1 -373
box -9 -175 424 100
use buff  buff_0
timestamp 1619185680
transform 1 0 446 0 1 -324
box 0 -49 54 51
use dff  dff_4
timestamp 1619465570
transform 1 0 587 0 1 -361
box 0 -201 239 89
<< labels >>
rlabel space 497 -328 497 -328 1 dc4
rlabel metal1 -184 630 -179 634 1 da1
rlabel metal1 119 630 124 634 1 da2
rlabel metal1 415 630 420 634 1 da3
rlabel metal1 727 630 732 634 1 da4
rlabel metal1 727 314 732 318 1 db4
rlabel metal1 415 314 420 318 1 db3
rlabel metal1 119 314 124 318 1 db2
rlabel metal1 -184 314 -179 318 1 db1
rlabel metal1 -65 -687 -60 -682 1 s1
rlabel metal1 -65 -796 -60 -791 1 s1_b
rlabel metal1 238 -796 243 -791 1 s2_b
rlabel metal1 238 -687 243 -682 1 s2
rlabel metal1 534 -687 539 -682 1 s3
rlabel metal1 534 -796 539 -791 1 s3_b
rlabel metal1 846 -796 851 -791 7 s4_b
rlabel metal1 846 -687 851 -682 7 s4
rlabel metal1 -350 675 -348 680 1 clk
rlabel metal1 361 71 364 72 1 gnd
rlabel metal1 821 -419 826 -415 1 c4_b
rlabel metal1 821 -307 826 -303 1 c4
rlabel metal1 115 -505 117 -502 1 ds1
rlabel metal1 217 -505 219 -502 1 ds2
rlabel metal1 318 -505 320 -502 1 ds3
rlabel m123contact 419 -506 424 -501 1 ds4
rlabel metal1 342 168 347 170 1 vdd
<< end >>
