magic
tech scmos
timestamp 1619185653
<< ntransistor >>
rect 11 12 13 17
rect 11 -23 13 -18
<< ndiffusion >>
rect 10 12 11 17
rect 13 12 14 17
rect 10 -23 11 -18
rect 13 -23 14 -18
<< ndcontact >>
rect 6 12 10 17
rect 14 12 18 17
rect 6 -23 10 -18
rect 14 -23 18 -18
<< polysilicon >>
rect 11 17 13 20
rect 11 -1 13 12
rect 11 -18 13 -6
rect 11 -26 13 -23
<< polycontact >>
rect 13 -1 17 4
rect 13 -13 17 -8
<< metal1 >>
rect 18 12 24 17
rect 6 -2 10 12
rect 17 -1 24 4
rect 3 -7 10 -2
rect 6 -18 10 -7
rect 17 -13 24 -8
rect 14 -27 18 -23
rect 0 -30 24 -27
<< end >>
