* SPICE3 file created from or.ext - technology: scmos

.option scale=0.09u

M1000 a_13_n29# a_11_n32# a_6_n29# Gnd nfet w=5 l=2
+  ad=25 pd=20 as=50 ps=40
M1001 a_13_8# a_11_n2# a_6_n29# Gnd nfet w=5 l=2
+  ad=25 pd=20 as=0 ps=0
