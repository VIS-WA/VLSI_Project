* SPICE3 file created from inv.ext - technology: scmos
Prop and Generate
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={5*LAMBDA}
.param width_P={10*LAMBDA}
.global gnd vdd

Vdd vdd gnd 'SUPPLY'
va1 in 0 pulse 0 1.8 0ns 0ns 0ns 10ns 20ns
va b 0 pulse 0 1.8 0ns 0ns 0ns 20ns 40ns
vb1 b_b 0 pulse 1.8 0 0ns 0ns 0ns 20ns 40ns
vb a_b 0 pulse 1.8 0 0ns 0ns 0ns 10ns 20ns

.option scale=0.09u

M1000 out in gnd Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=25 ps=20
M1001 out in vdd w_0_0# CMOSP w=10 l=2
+  ad=50 pd=30 as=50 ps=30
C0 in w_0_0# 0.08fF
C1 w_0_0# vdd 0.03fF
C2 in out 0.05fF
C3 out vdd 0.10fF
C4 w_0_0# out 0.04fF
C5 in gnd 0.05fF
C6 out gnd 0.05fF
C7 gnd Gnd 0.16fF
C8 out Gnd 0.04fF
C9 vdd Gnd 0.13fF
C10 in Gnd 0.14fF
C11 w_0_0# Gnd 0.58fF
.tran 0.1n 50n

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7)
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7)


run
plot v(in) v(out)



*hardcopy fig_inv_trans.eps v(b) v(c)
.endc

