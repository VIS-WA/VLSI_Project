4 bit CLA
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={5*LAMBDA}
.param width_P={10*LAMBDA}
.global gnd vdd

Vdd vdd gnd 'SUPPLY'


vp1 p1 0 pulse 1.8 1.8 0ns 1ns 1ns 10ns 20ns
vp2 p2 0 pulse 0 0 0ns 1ns 1ns 10ns 20ns
vp3 p3 0 pulse 0 0 0ns 1ns 1ns 10ns 20ns
vp4 p4 0 pulse 0 0 0ns 1ns 1ns 10ns 20ns

Vg1 g1 0 pulse 1.8 1.8 0ns 1ns 1ns 10ns 20ns $ select inv inputs
Vg2 g2 0 pulse 0 0 0ns 1ns 1ns 10ns 20ns $ select inv inputs
Vg3 g3 0 pulse 0 0 0ns 1ns 1ns 10ns 20ns $ select inv inputs
Vg4 g4 0 pulse 0 0 0ns 1ns 1ns 10ns 20ns $ select inv inputs

.option scale=0.09u

M1000 g4 z53 z54 Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=75 ps=60
M1001 vdd z53_b z54 Gnd CMOSN w=5 l=2
+  ad=175 pd=140 as=0 ps=0
M1002 z43 z41_b c3 Gnd CMOSN w=5 l=2
+  ad=75 pd=60 as=50 ps=40
M1003 vdd z41 c3 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 z54 m1_475_31# z55 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=75 ps=60
M1005 vdd m1_586_26# z55 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 z55 z51_b cc4 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=50 ps=40
M1007 vdd z51 cc4 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 g1_b g1 gnd Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=400 ps=320
M1009 g1_b g1 vdd vdd CMOSP w=10 l=2
+  ad=50 pd=30 as=450 ps=270
M1010 g2_b g2 gnd Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1011 g2_b g2 vdd vdd CMOSP w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1012 p3_b p3 gnd Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1013 p3_b p3 vdd vdd CMOSP w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1014 z41_b z41 gnd Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1015 z41_b z41 vdd vdd CMOSP w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1016 g3_b g3 gnd Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1017 g3_b g3 vdd vdd CMOSP w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1018 p4_b p4 gnd Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1019 p4_b p4 vdd vdd CMOSP w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1020 m1_586_26# m1_475_31# gnd Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1021 m1_586_26# m1_475_31# vdd vdd CMOSP w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1022 gnd g1_b c1 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=50 ps=40
M1023 vdd g1 c1 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 z51_b z51 gnd Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1025 z51_b z51 vdd vdd CMOSP w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1026 gnd g2 z42 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=75 ps=60
M1027 p3 g2_b z42 Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1028 z53_b z53 gnd Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1029 z53_b z53 vdd vdd CMOSP w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1030 gnd g1_b z2 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=100 ps=80
M1031 p2 g1 z2 Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1032 gnd p3_b z41 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=100 ps=80
M1033 z2 p3 z41 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 gnd p4_b m1_475_31# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=50 ps=40
M1035 z42 p4 m1_475_31# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 gnd p4_b z51 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=50 ps=40
M1037 z41 p4 z51 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 gnd p4_b z53 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=50 ps=40
M1039 g3 p4 z53 Gnd CMOSN w=5 l=2
+  ad=25 pd=20 as=0 ps=0
M1040 z2 g2_b c2 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=50 ps=40
M1041 vdd g2 c2 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 z41 g3_b z43 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 vdd g3 z43 Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd Gnd 6.50fF

.tran 0.1n 20n

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7)
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7)


run
plot v(c1) v(vdd) 
plot v(c2) v(vdd) 
plot v(c3) v(vdd) 
plot v(cc4) v(vdd) 
.endc
